#! /usr/bin/vvp
:ivl_version "12.0 (stable)";
:ivl_delay_selection "TYPICAL";
:vpi_time_precision + 0;
:vpi_module "/usr/lib/x86_64-linux-gnu/ivl/system.vpi";
:vpi_module "/usr/lib/x86_64-linux-gnu/ivl/vhdl_sys.vpi";
:vpi_module "/usr/lib/x86_64-linux-gnu/ivl/vhdl_textio.vpi";
:vpi_module "/usr/lib/x86_64-linux-gnu/ivl/v2005_math.vpi";
:vpi_module "/usr/lib/x86_64-linux-gnu/ivl/va_math.vpi";
S_0x5c7c329f9ad0 .scope module, "Add16" "Add16" 2 1;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "a";
    .port_info 1 /INPUT 16 "b";
    .port_info 2 /OUTPUT 16 "sum";
o0x7d2eeb85fac8 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c32f04ad0_0 .net "a", 15 0, o0x7d2eeb85fac8;  0 drivers
o0x7d2eeb85faf8 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c32f04bd0_0 .net "b", 15 0, o0x7d2eeb85faf8;  0 drivers
v0x5c7c32f04cb0_0 .net "c0", 0 0, L_0x5c7c33111ce0;  1 drivers
v0x5c7c32f04d50_0 .net "c1", 0 0, L_0x5c7c33114e80;  1 drivers
v0x5c7c32f04df0_0 .net "c10", 0 0, L_0x5c7c3312a3c0;  1 drivers
v0x5c7c32f04e90_0 .net "c11", 0 0, L_0x5c7c3312c930;  1 drivers
v0x5c7c32f04f30_0 .net "c12", 0 0, L_0x5c7c3312ef50;  1 drivers
v0x5c7c32f04fd0_0 .net "c13", 0 0, L_0x5c7c33131580;  1 drivers
v0x5c7c32f05070_0 .net "c14", 0 0, L_0x5c7c33133bc0;  1 drivers
v0x5c7c32f05110_0 .net "c15", 0 0, L_0x5c7c33136210;  1 drivers
v0x5c7c32f05240_0 .net "c2", 0 0, L_0x5c7c33117480;  1 drivers
v0x5c7c32f052e0_0 .net "c3", 0 0, L_0x5c7c33119a20;  1 drivers
v0x5c7c32f05380_0 .net "c4", 0 0, L_0x5c7c3311c0e0;  1 drivers
v0x5c7c32f05420_0 .net "c5", 0 0, L_0x5c7c3311e6a0;  1 drivers
v0x5c7c32f054c0_0 .net "c6", 0 0, L_0x5c7c33120bf0;  1 drivers
v0x5c7c32f05560_0 .net "c7", 0 0, L_0x5c7c33123160;  1 drivers
v0x5c7c32f05600_0 .net "c8", 0 0, L_0x5c7c33125850;  1 drivers
v0x5c7c32f057b0_0 .net "c9", 0 0, L_0x5c7c33127dc0;  1 drivers
v0x5c7c32f05850_0 .net "sum", 15 0, L_0x5c7c33136a20;  1 drivers
L_0x5c7c33112b10 .part o0x7d2eeb85fac8, 0, 1;
L_0x5c7c33112be0 .part o0x7d2eeb85faf8, 0, 1;
L_0x5c7c33115020 .part o0x7d2eeb85fac8, 1, 1;
L_0x5c7c331150c0 .part o0x7d2eeb85faf8, 1, 1;
L_0x5c7c33117620 .part o0x7d2eeb85fac8, 2, 1;
L_0x5c7c331176c0 .part o0x7d2eeb85faf8, 2, 1;
L_0x5c7c33119bc0 .part o0x7d2eeb85fac8, 3, 1;
L_0x5c7c33119c60 .part o0x7d2eeb85faf8, 3, 1;
L_0x5c7c3311c280 .part o0x7d2eeb85fac8, 4, 1;
L_0x5c7c3311c320 .part o0x7d2eeb85faf8, 4, 1;
L_0x5c7c3311e840 .part o0x7d2eeb85fac8, 5, 1;
L_0x5c7c3311e8e0 .part o0x7d2eeb85faf8, 5, 1;
L_0x5c7c33120d90 .part o0x7d2eeb85fac8, 6, 1;
L_0x5c7c33120e30 .part o0x7d2eeb85faf8, 6, 1;
L_0x5c7c33123300 .part o0x7d2eeb85fac8, 7, 1;
L_0x5c7c331234b0 .part o0x7d2eeb85faf8, 7, 1;
L_0x5c7c331259f0 .part o0x7d2eeb85fac8, 8, 1;
L_0x5c7c33125a90 .part o0x7d2eeb85faf8, 8, 1;
L_0x5c7c33127f60 .part o0x7d2eeb85fac8, 9, 1;
L_0x5c7c33128000 .part o0x7d2eeb85faf8, 9, 1;
L_0x5c7c33125b30 .part o0x7d2eeb85fac8, 10, 1;
L_0x5c7c3312a560 .part o0x7d2eeb85faf8, 10, 1;
L_0x5c7c3312cad0 .part o0x7d2eeb85fac8, 11, 1;
L_0x5c7c3312cb70 .part o0x7d2eeb85faf8, 11, 1;
L_0x5c7c3312f0f0 .part o0x7d2eeb85fac8, 12, 1;
L_0x5c7c3312f190 .part o0x7d2eeb85faf8, 12, 1;
L_0x5c7c33131720 .part o0x7d2eeb85fac8, 13, 1;
L_0x5c7c331317c0 .part o0x7d2eeb85faf8, 13, 1;
L_0x5c7c33133d60 .part o0x7d2eeb85fac8, 14, 1;
L_0x5c7c33133e00 .part o0x7d2eeb85faf8, 14, 1;
L_0x5c7c331363b0 .part o0x7d2eeb85fac8, 15, 1;
L_0x5c7c33136660 .part o0x7d2eeb85faf8, 15, 1;
LS_0x5c7c33136a20_0_0 .concat8 [ 1 1 1 1], L_0x5c7c33112950, L_0x5c7c331146d0, L_0x5c7c33116cd0, L_0x5c7c33119270;
LS_0x5c7c33136a20_0_4 .concat8 [ 1 1 1 1], L_0x5c7c3311b930, L_0x5c7c3311def0, L_0x5c7c33120440, L_0x5c7c331229b0;
LS_0x5c7c33136a20_0_8 .concat8 [ 1 1 1 1], L_0x5c7c331250a0, L_0x5c7c33127610, L_0x5c7c33129c10, L_0x5c7c3312c180;
LS_0x5c7c33136a20_0_12 .concat8 [ 1 1 1 1], L_0x5c7c3312e7a0, L_0x5c7c33130dd0, L_0x5c7c33133410, L_0x5c7c33135a60;
L_0x5c7c33136a20 .concat8 [ 4 4 4 4], LS_0x5c7c33136a20_0_0, LS_0x5c7c33136a20_0_4, LS_0x5c7c33136a20_0_8, LS_0x5c7c33136a20_0_12;
S_0x5c7c32d066a0 .scope module, "fa_gate10" "FullAdder" 2 15, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32d2c300_0 .net "a", 0 0, L_0x5c7c33127f60;  1 drivers
v0x5c7c32d2c3a0_0 .net "b", 0 0, L_0x5c7c33128000;  1 drivers
v0x5c7c32d2c460_0 .net "c", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d2c500_0 .net "carry", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d2c5a0_0 .net "sum", 0 0, L_0x5c7c33127610;  1 drivers
v0x5c7c32d2c640_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33125bd0;  1 drivers
v0x5c7c32d2c6e0_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33126ce0;  1 drivers
v0x5c7c32d2c780_0 .net "tmp_sum_out", 0 0, L_0x5c7c331266e0;  1 drivers
S_0x5c7c32d09150 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32d066a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d19ce0_0 .net "a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c8cd90_0 .net "b", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32d19fc0_0 .net "carry", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32d1a060_0 .net "sum", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
S_0x5c7c32d0bc00 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d09150;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32c7d6c0_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c94520_0 .net "in_b", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32c94140_0 .net "out", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32c893c0_0 .net "temp_out", 0 0, L_0x5c7c32ef7a00;  1 drivers
S_0x5c7c32d13c10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d0bc00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ef7a00 .functor NAND 1, L_0x5c7c33127f60, L_0x5c7c33128000, C4<1>, C4<1>;
v0x5c7c32cf67a0_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32cf3cf0_0 .net "in_b", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32cf1240_0 .net "out", 0 0, L_0x5c7c32ef7a00;  alias, 1 drivers
S_0x5c7c32d166c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d0bc00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32c7da50_0 .net "in_a", 0 0, L_0x5c7c32ef7a00;  alias, 1 drivers
v0x5c7c32c7db10_0 .net "out", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
S_0x5c7c32c7bec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d166c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125bd0 .functor NAND 1, L_0x5c7c32ef7a00, L_0x5c7c32ef7a00, C4<1>, C4<1>;
v0x5c7c32cee730_0 .net "in_a", 0 0, L_0x5c7c32ef7a00;  alias, 1 drivers
v0x5c7c32c7e6c0_0 .net "in_b", 0 0, L_0x5c7c32ef7a00;  alias, 1 drivers
v0x5c7c32c7e270_0 .net "out", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
S_0x5c7c32cc1b90 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d09150;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d19600_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32d196a0_0 .net "in_b", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32d19760_0 .net "out", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d19800_0 .net "temp_a_and_out", 0 0, L_0x5c7c33125da0;  1 drivers
v0x5c7c32d199b0_0 .net "temp_a_out", 0 0, L_0x5c7c33125c40;  1 drivers
v0x5c7c32d19a50_0 .net "temp_b_and_out", 0 0, L_0x5c7c33125fb0;  1 drivers
v0x5c7c32d19c00_0 .net "temp_b_out", 0 0, L_0x5c7c33125e50;  1 drivers
S_0x5c7c32cec350 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32cc1b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32c91a70_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c91b10_0 .net "in_b", 0 0, L_0x5c7c33125c40;  alias, 1 drivers
v0x5c7c32c890d0_0 .net "out", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
v0x5c7c32c91160_0 .net "temp_out", 0 0, L_0x5c7c33125cf0;  1 drivers
S_0x5c7c32c7c530 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32cec350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125cf0 .functor NAND 1, L_0x5c7c33127f60, L_0x5c7c33125c40, C4<1>, C4<1>;
v0x5c7c32c89460_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c93830_0 .net "in_b", 0 0, L_0x5c7c33125c40;  alias, 1 drivers
v0x5c7c32c938f0_0 .net "out", 0 0, L_0x5c7c33125cf0;  alias, 1 drivers
S_0x5c7c324ea9b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32cec350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32c91e50_0 .net "in_a", 0 0, L_0x5c7c33125cf0;  alias, 1 drivers
v0x5c7c32c91ef0_0 .net "out", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
S_0x5c7c324eab90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c324ea9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125da0 .functor NAND 1, L_0x5c7c33125cf0, L_0x5c7c33125cf0, C4<1>, C4<1>;
v0x5c7c32c93470_0 .net "in_a", 0 0, L_0x5c7c33125cf0;  alias, 1 drivers
v0x5c7c32c92b40_0 .net "in_b", 0 0, L_0x5c7c33125cf0;  alias, 1 drivers
v0x5c7c32c92760_0 .net "out", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
S_0x5c7c324ebdc0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32cc1b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32c8f3a0_0 .net "in_a", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32c8f440_0 .net "in_b", 0 0, L_0x5c7c33125e50;  alias, 1 drivers
v0x5c7c32c8ea90_0 .net "out", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
v0x5c7c32c8e6b0_0 .net "temp_out", 0 0, L_0x5c7c33125f00;  1 drivers
S_0x5c7c324ebfa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c324ebdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125f00 .functor NAND 1, L_0x5c7c33128000, L_0x5c7c33125e50, C4<1>, C4<1>;
v0x5c7c32c91220_0 .net "in_a", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32c90d80_0 .net "in_b", 0 0, L_0x5c7c33125e50;  alias, 1 drivers
v0x5c7c32c90e40_0 .net "out", 0 0, L_0x5c7c33125f00;  alias, 1 drivers
S_0x5c7c324d2890 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c324ebdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32c8f780_0 .net "in_a", 0 0, L_0x5c7c33125f00;  alias, 1 drivers
v0x5c7c32c8f820_0 .net "out", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
S_0x5c7c324d2a70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c324d2890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125fb0 .functor NAND 1, L_0x5c7c33125f00, L_0x5c7c33125f00, C4<1>, C4<1>;
v0x5c7c32c90470_0 .net "in_a", 0 0, L_0x5c7c33125f00;  alias, 1 drivers
v0x5c7c32c90530_0 .net "in_b", 0 0, L_0x5c7c33125f00;  alias, 1 drivers
v0x5c7c32c900e0_0 .net "out", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
S_0x5c7c324d42f0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32cc1b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32c8d0b0_0 .net "in_a", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32c8d150_0 .net "out", 0 0, L_0x5c7c33125c40;  alias, 1 drivers
S_0x5c7c324d4480 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c324d42f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125c40 .functor NAND 1, L_0x5c7c33128000, L_0x5c7c33128000, C4<1>, C4<1>;
v0x5c7c324d46d0_0 .net "in_a", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32c8de30_0 .net "in_b", 0 0, L_0x5c7c33128000;  alias, 1 drivers
v0x5c7c32c8d9c0_0 .net "out", 0 0, L_0x5c7c33125c40;  alias, 1 drivers
S_0x5c7c324c9360 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32cc1b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32c8c070_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c88a60_0 .net "out", 0 0, L_0x5c7c33125e50;  alias, 1 drivers
S_0x5c7c324c9540 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c324c9360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125e50 .functor NAND 1, L_0x5c7c33127f60, L_0x5c7c33127f60, C4<1>, C4<1>;
v0x5c7c32c8ccd0_0 .net "in_a", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c8c3c0_0 .net "in_b", 0 0, L_0x5c7c33127f60;  alias, 1 drivers
v0x5c7c32c8c480_0 .net "out", 0 0, L_0x5c7c33125e50;  alias, 1 drivers
S_0x5c7c324d6930 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32cc1b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d18f50_0 .net "branch1_out", 0 0, L_0x5c7c331261c0;  1 drivers
v0x5c7c32d19080_0 .net "branch2_out", 0 0, L_0x5c7c33126450;  1 drivers
v0x5c7c32d191d0_0 .net "in_a", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
v0x5c7c32d192a0_0 .net "in_b", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
v0x5c7c32d19340_0 .net "out", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d193e0_0 .net "temp1_out", 0 0, L_0x5c7c33126110;  1 drivers
v0x5c7c32d19480_0 .net "temp2_out", 0 0, L_0x5c7c331263a0;  1 drivers
v0x5c7c32d19520_0 .net "temp3_out", 0 0, L_0x5c7c33126630;  1 drivers
S_0x5c7c324d6bb0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c324d6930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32c89aa0_0 .net "in_a", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
v0x5c7c32c89b40_0 .net "in_b", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
v0x5c7c32c92110_0 .net "out", 0 0, L_0x5c7c33126110;  alias, 1 drivers
v0x5c7c32c60d10_0 .net "temp_out", 0 0, L_0x5c7c33126060;  1 drivers
S_0x5c7c324e8930 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c324d6bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126060 .functor NAND 1, L_0x5c7c33125da0, L_0x5c7c33125da0, C4<1>, C4<1>;
v0x5c7c324e8b60_0 .net "in_a", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
v0x5c7c324e8c20_0 .net "in_b", 0 0, L_0x5c7c33125da0;  alias, 1 drivers
v0x5c7c32c8b6d0_0 .net "out", 0 0, L_0x5c7c33126060;  alias, 1 drivers
S_0x5c7c324f3080 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c324d6bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32c89e30_0 .net "in_a", 0 0, L_0x5c7c33126060;  alias, 1 drivers
v0x5c7c32c89ed0_0 .net "out", 0 0, L_0x5c7c33126110;  alias, 1 drivers
S_0x5c7c324f3210 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c324f3080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126110 .functor NAND 1, L_0x5c7c33126060, L_0x5c7c33126060, C4<1>, C4<1>;
v0x5c7c32c8b2f0_0 .net "in_a", 0 0, L_0x5c7c33126060;  alias, 1 drivers
v0x5c7c32c8a9e0_0 .net "in_b", 0 0, L_0x5c7c33126060;  alias, 1 drivers
v0x5c7c32c8a650_0 .net "out", 0 0, L_0x5c7c33126110;  alias, 1 drivers
S_0x5c7c324e5940 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c324d6930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c324cb4e0_0 .net "in_a", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
v0x5c7c324cb580_0 .net "in_b", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
v0x5c7c324cb620_0 .net "out", 0 0, L_0x5c7c331263a0;  alias, 1 drivers
v0x5c7c324cb740_0 .net "temp_out", 0 0, L_0x5c7c32d179d0;  1 drivers
S_0x5c7c324e5b20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c324e5940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d179d0 .functor NAND 1, L_0x5c7c33125fb0, L_0x5c7c33125fb0, C4<1>, C4<1>;
v0x5c7c32c836b0_0 .net "in_a", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
v0x5c7c32c83770_0 .net "in_b", 0 0, L_0x5c7c33125fb0;  alias, 1 drivers
v0x5c7c32ce9510_0 .net "out", 0 0, L_0x5c7c32d179d0;  alias, 1 drivers
S_0x5c7c32490490 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c324e5940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c324d1dd0_0 .net "in_a", 0 0, L_0x5c7c32d179d0;  alias, 1 drivers
v0x5c7c324d1e70_0 .net "out", 0 0, L_0x5c7c331263a0;  alias, 1 drivers
S_0x5c7c32490620 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32490490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331263a0 .functor NAND 1, L_0x5c7c32d179d0, L_0x5c7c32d179d0, C4<1>, C4<1>;
v0x5c7c324d1b20_0 .net "in_a", 0 0, L_0x5c7c32d179d0;  alias, 1 drivers
v0x5c7c324d1be0_0 .net "in_b", 0 0, L_0x5c7c32d179d0;  alias, 1 drivers
v0x5c7c324d1cd0_0 .net "out", 0 0, L_0x5c7c331263a0;  alias, 1 drivers
S_0x5c7c324e3330 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c324d6930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d171d0_0 .net "in_a", 0 0, L_0x5c7c331261c0;  alias, 1 drivers
v0x5c7c32d17270_0 .net "in_b", 0 0, L_0x5c7c33126450;  alias, 1 drivers
v0x5c7c32d17310_0 .net "out", 0 0, L_0x5c7c33126630;  alias, 1 drivers
v0x5c7c32d173b0_0 .net "temp_out", 0 0, L_0x5c7c32d18340;  1 drivers
S_0x5c7c324e3510 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c324e3330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d18340 .functor NAND 1, L_0x5c7c331261c0, L_0x5c7c33126450, C4<1>, C4<1>;
v0x5c7c324cb8b0_0 .net "in_a", 0 0, L_0x5c7c331261c0;  alias, 1 drivers
v0x5c7c324d7eb0_0 .net "in_b", 0 0, L_0x5c7c33126450;  alias, 1 drivers
v0x5c7c324d7f70_0 .net "out", 0 0, L_0x5c7c32d18340;  alias, 1 drivers
S_0x5c7c324d80c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c324e3330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d17090_0 .net "in_a", 0 0, L_0x5c7c32d18340;  alias, 1 drivers
v0x5c7c32d17130_0 .net "out", 0 0, L_0x5c7c33126630;  alias, 1 drivers
S_0x5c7c324da150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c324d80c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126630 .functor NAND 1, L_0x5c7c32d18340, L_0x5c7c32d18340, C4<1>, C4<1>;
v0x5c7c324da370_0 .net "in_a", 0 0, L_0x5c7c32d18340;  alias, 1 drivers
v0x5c7c324da460_0 .net "in_b", 0 0, L_0x5c7c32d18340;  alias, 1 drivers
v0x5c7c32d16ff0_0 .net "out", 0 0, L_0x5c7c33126630;  alias, 1 drivers
S_0x5c7c32d174e0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c324d6930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d17b20_0 .net "in_a", 0 0, L_0x5c7c33126110;  alias, 1 drivers
v0x5c7c32d17bc0_0 .net "out", 0 0, L_0x5c7c331261c0;  alias, 1 drivers
S_0x5c7c32d17670 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d174e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331261c0 .functor NAND 1, L_0x5c7c33126110, L_0x5c7c33126110, C4<1>, C4<1>;
v0x5c7c32d17850_0 .net "in_a", 0 0, L_0x5c7c33126110;  alias, 1 drivers
v0x5c7c32d178f0_0 .net "in_b", 0 0, L_0x5c7c33126110;  alias, 1 drivers
v0x5c7c32d17a40_0 .net "out", 0 0, L_0x5c7c331261c0;  alias, 1 drivers
S_0x5c7c32d17cc0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c324d6930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d18490_0 .net "in_a", 0 0, L_0x5c7c331263a0;  alias, 1 drivers
v0x5c7c32d18530_0 .net "out", 0 0, L_0x5c7c33126450;  alias, 1 drivers
S_0x5c7c32d17f30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d17cc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126450 .functor NAND 1, L_0x5c7c331263a0, L_0x5c7c331263a0, C4<1>, C4<1>;
v0x5c7c32d181a0_0 .net "in_a", 0 0, L_0x5c7c331263a0;  alias, 1 drivers
v0x5c7c32d18260_0 .net "in_b", 0 0, L_0x5c7c331263a0;  alias, 1 drivers
v0x5c7c32d183b0_0 .net "out", 0 0, L_0x5c7c33126450;  alias, 1 drivers
S_0x5c7c32d18630 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c324d6930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d18dd0_0 .net "in_a", 0 0, L_0x5c7c33126630;  alias, 1 drivers
v0x5c7c32d18e70_0 .net "out", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
S_0x5c7c32d18850 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d18630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331266e0 .functor NAND 1, L_0x5c7c33126630, L_0x5c7c33126630, C4<1>, C4<1>;
v0x5c7c32d18ac0_0 .net "in_a", 0 0, L_0x5c7c33126630;  alias, 1 drivers
v0x5c7c32d18b80_0 .net "in_b", 0 0, L_0x5c7c33126630;  alias, 1 drivers
v0x5c7c32d18cd0_0 .net "out", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
S_0x5c7c32d1a140 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32d066a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d25c50_0 .net "a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d25cf0_0 .net "b", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d25ec0_0 .net "carry", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d25f60_0 .net "sum", 0 0, L_0x5c7c33127610;  alias, 1 drivers
S_0x5c7c32d1a2f0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d1a140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d1b300_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1b3a0_0 .net "in_b", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1b490_0 .net "out", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d1b5b0_0 .net "temp_out", 0 0, L_0x5c7c32d18c60;  1 drivers
S_0x5c7c32d1a4a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d1a2f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d18c60 .functor NAND 1, L_0x5c7c331266e0, L_0x5c7c33125850, C4<1>, C4<1>;
v0x5c7c32d1a710_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1a7d0_0 .net "in_b", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1a890_0 .net "out", 0 0, L_0x5c7c32d18c60;  alias, 1 drivers
S_0x5c7c32d1a9e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d1a2f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d1b150_0 .net "in_a", 0 0, L_0x5c7c32d18c60;  alias, 1 drivers
v0x5c7c32d1b1f0_0 .net "out", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
S_0x5c7c32d1ac00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d1a9e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126ce0 .functor NAND 1, L_0x5c7c32d18c60, L_0x5c7c32d18c60, C4<1>, C4<1>;
v0x5c7c32d1ae70_0 .net "in_a", 0 0, L_0x5c7c32d18c60;  alias, 1 drivers
v0x5c7c32d1af60_0 .net "in_b", 0 0, L_0x5c7c32d18c60;  alias, 1 drivers
v0x5c7c32d1b050_0 .net "out", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
S_0x5c7c32d1b700 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d1a140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d25570_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d25610_0 .net "in_b", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d256d0_0 .net "out", 0 0, L_0x5c7c33127610;  alias, 1 drivers
v0x5c7c32d25770_0 .net "temp_a_and_out", 0 0, L_0x5c7c33126ef0;  1 drivers
v0x5c7c32d25920_0 .net "temp_a_out", 0 0, L_0x5c7c33126d90;  1 drivers
v0x5c7c32d259c0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33127100;  1 drivers
v0x5c7c32d25b70_0 .net "temp_b_out", 0 0, L_0x5c7c33126fa0;  1 drivers
S_0x5c7c32d1b8e0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d1b700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d1c980_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1cb30_0 .net "in_b", 0 0, L_0x5c7c33126d90;  alias, 1 drivers
v0x5c7c32d1cc20_0 .net "out", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
v0x5c7c32d1cd40_0 .net "temp_out", 0 0, L_0x5c7c33126e40;  1 drivers
S_0x5c7c32d1bb50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d1b8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126e40 .functor NAND 1, L_0x5c7c331266e0, L_0x5c7c33126d90, C4<1>, C4<1>;
v0x5c7c32d1bdc0_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1be80_0 .net "in_b", 0 0, L_0x5c7c33126d90;  alias, 1 drivers
v0x5c7c32d1bf40_0 .net "out", 0 0, L_0x5c7c33126e40;  alias, 1 drivers
S_0x5c7c32d1c060 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d1b8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d1c7d0_0 .net "in_a", 0 0, L_0x5c7c33126e40;  alias, 1 drivers
v0x5c7c32d1c870_0 .net "out", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
S_0x5c7c32d1c280 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d1c060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126ef0 .functor NAND 1, L_0x5c7c33126e40, L_0x5c7c33126e40, C4<1>, C4<1>;
v0x5c7c32d1c4f0_0 .net "in_a", 0 0, L_0x5c7c33126e40;  alias, 1 drivers
v0x5c7c32d1c5e0_0 .net "in_b", 0 0, L_0x5c7c33126e40;  alias, 1 drivers
v0x5c7c32d1c6d0_0 .net "out", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
S_0x5c7c32d1ce00 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d1b700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d1de30_0 .net "in_a", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1ded0_0 .net "in_b", 0 0, L_0x5c7c33126fa0;  alias, 1 drivers
v0x5c7c32d1dfc0_0 .net "out", 0 0, L_0x5c7c33127100;  alias, 1 drivers
v0x5c7c32d1e0e0_0 .net "temp_out", 0 0, L_0x5c7c33127050;  1 drivers
S_0x5c7c32d1cfe0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d1ce00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127050 .functor NAND 1, L_0x5c7c33125850, L_0x5c7c33126fa0, C4<1>, C4<1>;
v0x5c7c32d1d250_0 .net "in_a", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1d360_0 .net "in_b", 0 0, L_0x5c7c33126fa0;  alias, 1 drivers
v0x5c7c32d1d420_0 .net "out", 0 0, L_0x5c7c33127050;  alias, 1 drivers
S_0x5c7c32d1d540 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d1ce00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d1dc80_0 .net "in_a", 0 0, L_0x5c7c33127050;  alias, 1 drivers
v0x5c7c32d1dd20_0 .net "out", 0 0, L_0x5c7c33127100;  alias, 1 drivers
S_0x5c7c32d1d760 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d1d540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127100 .functor NAND 1, L_0x5c7c33127050, L_0x5c7c33127050, C4<1>, C4<1>;
v0x5c7c32d1d9d0_0 .net "in_a", 0 0, L_0x5c7c33127050;  alias, 1 drivers
v0x5c7c32d1da90_0 .net "in_b", 0 0, L_0x5c7c33127050;  alias, 1 drivers
v0x5c7c32d1db80_0 .net "out", 0 0, L_0x5c7c33127100;  alias, 1 drivers
S_0x5c7c32d1e230 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d1b700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d1e970_0 .net "in_a", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1ea10_0 .net "out", 0 0, L_0x5c7c33126d90;  alias, 1 drivers
S_0x5c7c32d1e400 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d1e230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126d90 .functor NAND 1, L_0x5c7c33125850, L_0x5c7c33125850, C4<1>, C4<1>;
v0x5c7c32d1e650_0 .net "in_a", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1e7a0_0 .net "in_b", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32d1e860_0 .net "out", 0 0, L_0x5c7c33126d90;  alias, 1 drivers
S_0x5c7c32d1eb10 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d1b700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d1f250_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1f2f0_0 .net "out", 0 0, L_0x5c7c33126fa0;  alias, 1 drivers
S_0x5c7c32d1ed30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d1eb10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33126fa0 .functor NAND 1, L_0x5c7c331266e0, L_0x5c7c331266e0, C4<1>, C4<1>;
v0x5c7c32d1efa0_0 .net "in_a", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1f060_0 .net "in_b", 0 0, L_0x5c7c331266e0;  alias, 1 drivers
v0x5c7c32d1f120_0 .net "out", 0 0, L_0x5c7c33126fa0;  alias, 1 drivers
S_0x5c7c32d1f3f0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d1b700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d24ec0_0 .net "branch1_out", 0 0, L_0x5c7c33127310;  1 drivers
v0x5c7c32d24ff0_0 .net "branch2_out", 0 0, L_0x5c7c33127490;  1 drivers
v0x5c7c32d25140_0 .net "in_a", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
v0x5c7c32d25210_0 .net "in_b", 0 0, L_0x5c7c33127100;  alias, 1 drivers
v0x5c7c32d252b0_0 .net "out", 0 0, L_0x5c7c33127610;  alias, 1 drivers
v0x5c7c32d25350_0 .net "temp1_out", 0 0, L_0x5c7c33127260;  1 drivers
v0x5c7c32d253f0_0 .net "temp2_out", 0 0, L_0x5c7c331273e0;  1 drivers
v0x5c7c32d25490_0 .net "temp3_out", 0 0, L_0x5c7c33127560;  1 drivers
S_0x5c7c32d1f670 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d1f3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d20700_0 .net "in_a", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
v0x5c7c32d207a0_0 .net "in_b", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
v0x5c7c32d20860_0 .net "out", 0 0, L_0x5c7c33127260;  alias, 1 drivers
v0x5c7c32d20980_0 .net "temp_out", 0 0, L_0x5c7c331271b0;  1 drivers
S_0x5c7c32d1f8e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d1f670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331271b0 .functor NAND 1, L_0x5c7c33126ef0, L_0x5c7c33126ef0, C4<1>, C4<1>;
v0x5c7c32d1fb50_0 .net "in_a", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
v0x5c7c32d1fc10_0 .net "in_b", 0 0, L_0x5c7c33126ef0;  alias, 1 drivers
v0x5c7c32d1fd60_0 .net "out", 0 0, L_0x5c7c331271b0;  alias, 1 drivers
S_0x5c7c32d1fe60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d1f670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d20550_0 .net "in_a", 0 0, L_0x5c7c331271b0;  alias, 1 drivers
v0x5c7c32d205f0_0 .net "out", 0 0, L_0x5c7c33127260;  alias, 1 drivers
S_0x5c7c32d20030 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d1fe60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127260 .functor NAND 1, L_0x5c7c331271b0, L_0x5c7c331271b0, C4<1>, C4<1>;
v0x5c7c32d202a0_0 .net "in_a", 0 0, L_0x5c7c331271b0;  alias, 1 drivers
v0x5c7c32d20360_0 .net "in_b", 0 0, L_0x5c7c331271b0;  alias, 1 drivers
v0x5c7c32d20450_0 .net "out", 0 0, L_0x5c7c33127260;  alias, 1 drivers
S_0x5c7c32d20af0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d1f3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d21b20_0 .net "in_a", 0 0, L_0x5c7c33127100;  alias, 1 drivers
v0x5c7c32d21bc0_0 .net "in_b", 0 0, L_0x5c7c33127100;  alias, 1 drivers
v0x5c7c32d21c80_0 .net "out", 0 0, L_0x5c7c331273e0;  alias, 1 drivers
v0x5c7c32d21da0_0 .net "temp_out", 0 0, L_0x5c7c32d23940;  1 drivers
S_0x5c7c32d20cd0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d20af0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d23940 .functor NAND 1, L_0x5c7c33127100, L_0x5c7c33127100, C4<1>, C4<1>;
v0x5c7c32d20f40_0 .net "in_a", 0 0, L_0x5c7c33127100;  alias, 1 drivers
v0x5c7c32d21000_0 .net "in_b", 0 0, L_0x5c7c33127100;  alias, 1 drivers
v0x5c7c32d21150_0 .net "out", 0 0, L_0x5c7c32d23940;  alias, 1 drivers
S_0x5c7c32d21250 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d20af0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d21970_0 .net "in_a", 0 0, L_0x5c7c32d23940;  alias, 1 drivers
v0x5c7c32d21a10_0 .net "out", 0 0, L_0x5c7c331273e0;  alias, 1 drivers
S_0x5c7c32d21420 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d21250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331273e0 .functor NAND 1, L_0x5c7c32d23940, L_0x5c7c32d23940, C4<1>, C4<1>;
v0x5c7c32d21690_0 .net "in_a", 0 0, L_0x5c7c32d23940;  alias, 1 drivers
v0x5c7c32d21780_0 .net "in_b", 0 0, L_0x5c7c32d23940;  alias, 1 drivers
v0x5c7c32d21870_0 .net "out", 0 0, L_0x5c7c331273e0;  alias, 1 drivers
S_0x5c7c32d21f10 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d1f3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d22f50_0 .net "in_a", 0 0, L_0x5c7c33127310;  alias, 1 drivers
v0x5c7c32d23020_0 .net "in_b", 0 0, L_0x5c7c33127490;  alias, 1 drivers
v0x5c7c32d230f0_0 .net "out", 0 0, L_0x5c7c33127560;  alias, 1 drivers
v0x5c7c32d23210_0 .net "temp_out", 0 0, L_0x5c7c32d242b0;  1 drivers
S_0x5c7c32d220f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d21f10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d242b0 .functor NAND 1, L_0x5c7c33127310, L_0x5c7c33127490, C4<1>, C4<1>;
v0x5c7c32d22340_0 .net "in_a", 0 0, L_0x5c7c33127310;  alias, 1 drivers
v0x5c7c32d22420_0 .net "in_b", 0 0, L_0x5c7c33127490;  alias, 1 drivers
v0x5c7c32d224e0_0 .net "out", 0 0, L_0x5c7c32d242b0;  alias, 1 drivers
S_0x5c7c32d22630 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d21f10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d22da0_0 .net "in_a", 0 0, L_0x5c7c32d242b0;  alias, 1 drivers
v0x5c7c32d22e40_0 .net "out", 0 0, L_0x5c7c33127560;  alias, 1 drivers
S_0x5c7c32d22850 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d22630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127560 .functor NAND 1, L_0x5c7c32d242b0, L_0x5c7c32d242b0, C4<1>, C4<1>;
v0x5c7c32d22ac0_0 .net "in_a", 0 0, L_0x5c7c32d242b0;  alias, 1 drivers
v0x5c7c32d22bb0_0 .net "in_b", 0 0, L_0x5c7c32d242b0;  alias, 1 drivers
v0x5c7c32d22ca0_0 .net "out", 0 0, L_0x5c7c33127560;  alias, 1 drivers
S_0x5c7c32d23360 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d1f3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d23a90_0 .net "in_a", 0 0, L_0x5c7c33127260;  alias, 1 drivers
v0x5c7c32d23b30_0 .net "out", 0 0, L_0x5c7c33127310;  alias, 1 drivers
S_0x5c7c32d23530 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d23360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127310 .functor NAND 1, L_0x5c7c33127260, L_0x5c7c33127260, C4<1>, C4<1>;
v0x5c7c32d237a0_0 .net "in_a", 0 0, L_0x5c7c33127260;  alias, 1 drivers
v0x5c7c32d23860_0 .net "in_b", 0 0, L_0x5c7c33127260;  alias, 1 drivers
v0x5c7c32d239b0_0 .net "out", 0 0, L_0x5c7c33127310;  alias, 1 drivers
S_0x5c7c32d23c30 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d1f3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d24400_0 .net "in_a", 0 0, L_0x5c7c331273e0;  alias, 1 drivers
v0x5c7c32d244a0_0 .net "out", 0 0, L_0x5c7c33127490;  alias, 1 drivers
S_0x5c7c32d23ea0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d23c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127490 .functor NAND 1, L_0x5c7c331273e0, L_0x5c7c331273e0, C4<1>, C4<1>;
v0x5c7c32d24110_0 .net "in_a", 0 0, L_0x5c7c331273e0;  alias, 1 drivers
v0x5c7c32d241d0_0 .net "in_b", 0 0, L_0x5c7c331273e0;  alias, 1 drivers
v0x5c7c32d24320_0 .net "out", 0 0, L_0x5c7c33127490;  alias, 1 drivers
S_0x5c7c32d245a0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d1f3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d24d40_0 .net "in_a", 0 0, L_0x5c7c33127560;  alias, 1 drivers
v0x5c7c32d24de0_0 .net "out", 0 0, L_0x5c7c33127610;  alias, 1 drivers
S_0x5c7c32d247c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d245a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127610 .functor NAND 1, L_0x5c7c33127560, L_0x5c7c33127560, C4<1>, C4<1>;
v0x5c7c32d24a30_0 .net "in_a", 0 0, L_0x5c7c33127560;  alias, 1 drivers
v0x5c7c32d24af0_0 .net "in_b", 0 0, L_0x5c7c33127560;  alias, 1 drivers
v0x5c7c32d24c40_0 .net "out", 0 0, L_0x5c7c33127610;  alias, 1 drivers
S_0x5c7c32d26040 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32d066a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d2ba30_0 .net "branch1_out", 0 0, L_0x5c7c331278a0;  1 drivers
v0x5c7c32d2bb60_0 .net "branch2_out", 0 0, L_0x5c7c33127b30;  1 drivers
v0x5c7c32d2bcb0_0 .net "in_a", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32d2be90_0 .net "in_b", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d2c040_0 .net "out", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d2c0e0_0 .net "temp1_out", 0 0, L_0x5c7c331277f0;  1 drivers
v0x5c7c32d2c180_0 .net "temp2_out", 0 0, L_0x5c7c33127a80;  1 drivers
v0x5c7c32d2c220_0 .net "temp3_out", 0 0, L_0x5c7c33127d10;  1 drivers
S_0x5c7c32d261d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d26040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d27270_0 .net "in_a", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32d27310_0 .net "in_b", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32d273d0_0 .net "out", 0 0, L_0x5c7c331277f0;  alias, 1 drivers
v0x5c7c32d274f0_0 .net "temp_out", 0 0, L_0x5c7c32d24bd0;  1 drivers
S_0x5c7c32d263f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d261d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d24bd0 .functor NAND 1, L_0x5c7c33125bd0, L_0x5c7c33125bd0, C4<1>, C4<1>;
v0x5c7c32d26660_0 .net "in_a", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32d267b0_0 .net "in_b", 0 0, L_0x5c7c33125bd0;  alias, 1 drivers
v0x5c7c32d26870_0 .net "out", 0 0, L_0x5c7c32d24bd0;  alias, 1 drivers
S_0x5c7c32d269a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d261d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d270c0_0 .net "in_a", 0 0, L_0x5c7c32d24bd0;  alias, 1 drivers
v0x5c7c32d27160_0 .net "out", 0 0, L_0x5c7c331277f0;  alias, 1 drivers
S_0x5c7c32d26b70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d269a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331277f0 .functor NAND 1, L_0x5c7c32d24bd0, L_0x5c7c32d24bd0, C4<1>, C4<1>;
v0x5c7c32d26de0_0 .net "in_a", 0 0, L_0x5c7c32d24bd0;  alias, 1 drivers
v0x5c7c32d26ed0_0 .net "in_b", 0 0, L_0x5c7c32d24bd0;  alias, 1 drivers
v0x5c7c32d26fc0_0 .net "out", 0 0, L_0x5c7c331277f0;  alias, 1 drivers
S_0x5c7c32d27660 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d26040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d28690_0 .net "in_a", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d28730_0 .net "in_b", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d287f0_0 .net "out", 0 0, L_0x5c7c33127a80;  alias, 1 drivers
v0x5c7c32d28910_0 .net "temp_out", 0 0, L_0x5c7c32d2a4b0;  1 drivers
S_0x5c7c32d27840 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d27660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d2a4b0 .functor NAND 1, L_0x5c7c33126ce0, L_0x5c7c33126ce0, C4<1>, C4<1>;
v0x5c7c32d27ab0_0 .net "in_a", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d27c00_0 .net "in_b", 0 0, L_0x5c7c33126ce0;  alias, 1 drivers
v0x5c7c32d27cc0_0 .net "out", 0 0, L_0x5c7c32d2a4b0;  alias, 1 drivers
S_0x5c7c32d27dc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d27660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d284e0_0 .net "in_a", 0 0, L_0x5c7c32d2a4b0;  alias, 1 drivers
v0x5c7c32d28580_0 .net "out", 0 0, L_0x5c7c33127a80;  alias, 1 drivers
S_0x5c7c32d27f90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d27dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127a80 .functor NAND 1, L_0x5c7c32d2a4b0, L_0x5c7c32d2a4b0, C4<1>, C4<1>;
v0x5c7c32d28200_0 .net "in_a", 0 0, L_0x5c7c32d2a4b0;  alias, 1 drivers
v0x5c7c32d282f0_0 .net "in_b", 0 0, L_0x5c7c32d2a4b0;  alias, 1 drivers
v0x5c7c32d283e0_0 .net "out", 0 0, L_0x5c7c33127a80;  alias, 1 drivers
S_0x5c7c32d28a80 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d26040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d29ac0_0 .net "in_a", 0 0, L_0x5c7c331278a0;  alias, 1 drivers
v0x5c7c32d29b90_0 .net "in_b", 0 0, L_0x5c7c33127b30;  alias, 1 drivers
v0x5c7c32d29c60_0 .net "out", 0 0, L_0x5c7c33127d10;  alias, 1 drivers
v0x5c7c32d29d80_0 .net "temp_out", 0 0, L_0x5c7c32d2ae20;  1 drivers
S_0x5c7c32d28c60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d28a80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d2ae20 .functor NAND 1, L_0x5c7c331278a0, L_0x5c7c33127b30, C4<1>, C4<1>;
v0x5c7c32d28eb0_0 .net "in_a", 0 0, L_0x5c7c331278a0;  alias, 1 drivers
v0x5c7c32d28f90_0 .net "in_b", 0 0, L_0x5c7c33127b30;  alias, 1 drivers
v0x5c7c32d29050_0 .net "out", 0 0, L_0x5c7c32d2ae20;  alias, 1 drivers
S_0x5c7c32d291a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d28a80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d29910_0 .net "in_a", 0 0, L_0x5c7c32d2ae20;  alias, 1 drivers
v0x5c7c32d299b0_0 .net "out", 0 0, L_0x5c7c33127d10;  alias, 1 drivers
S_0x5c7c32d293c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d291a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127d10 .functor NAND 1, L_0x5c7c32d2ae20, L_0x5c7c32d2ae20, C4<1>, C4<1>;
v0x5c7c32d29630_0 .net "in_a", 0 0, L_0x5c7c32d2ae20;  alias, 1 drivers
v0x5c7c32d29720_0 .net "in_b", 0 0, L_0x5c7c32d2ae20;  alias, 1 drivers
v0x5c7c32d29810_0 .net "out", 0 0, L_0x5c7c33127d10;  alias, 1 drivers
S_0x5c7c32d29ed0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d26040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d2a600_0 .net "in_a", 0 0, L_0x5c7c331277f0;  alias, 1 drivers
v0x5c7c32d2a6a0_0 .net "out", 0 0, L_0x5c7c331278a0;  alias, 1 drivers
S_0x5c7c32d2a0a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d29ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331278a0 .functor NAND 1, L_0x5c7c331277f0, L_0x5c7c331277f0, C4<1>, C4<1>;
v0x5c7c32d2a310_0 .net "in_a", 0 0, L_0x5c7c331277f0;  alias, 1 drivers
v0x5c7c32d2a3d0_0 .net "in_b", 0 0, L_0x5c7c331277f0;  alias, 1 drivers
v0x5c7c32d2a520_0 .net "out", 0 0, L_0x5c7c331278a0;  alias, 1 drivers
S_0x5c7c32d2a7a0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d26040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d2af70_0 .net "in_a", 0 0, L_0x5c7c33127a80;  alias, 1 drivers
v0x5c7c32d2b010_0 .net "out", 0 0, L_0x5c7c33127b30;  alias, 1 drivers
S_0x5c7c32d2aa10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d2a7a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127b30 .functor NAND 1, L_0x5c7c33127a80, L_0x5c7c33127a80, C4<1>, C4<1>;
v0x5c7c32d2ac80_0 .net "in_a", 0 0, L_0x5c7c33127a80;  alias, 1 drivers
v0x5c7c32d2ad40_0 .net "in_b", 0 0, L_0x5c7c33127a80;  alias, 1 drivers
v0x5c7c32d2ae90_0 .net "out", 0 0, L_0x5c7c33127b30;  alias, 1 drivers
S_0x5c7c32d2b110 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d26040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d2b8b0_0 .net "in_a", 0 0, L_0x5c7c33127d10;  alias, 1 drivers
v0x5c7c32d2b950_0 .net "out", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
S_0x5c7c32d2b330 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d2b110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33127dc0 .functor NAND 1, L_0x5c7c33127d10, L_0x5c7c33127d10, C4<1>, C4<1>;
v0x5c7c32d2b5a0_0 .net "in_a", 0 0, L_0x5c7c33127d10;  alias, 1 drivers
v0x5c7c32d2b660_0 .net "in_b", 0 0, L_0x5c7c33127d10;  alias, 1 drivers
v0x5c7c32d2b7b0_0 .net "out", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
S_0x5c7c32d2c880 .scope module, "fa_gate11" "FullAdder" 2 16, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32d4ab50_0 .net "a", 0 0, L_0x5c7c33125b30;  1 drivers
v0x5c7c32d4abf0_0 .net "b", 0 0, L_0x5c7c3312a560;  1 drivers
v0x5c7c32d4acb0_0 .net "c", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d4ad50_0 .net "carry", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d4adf0_0 .net "sum", 0 0, L_0x5c7c33129c10;  1 drivers
v0x5c7c32d4ae90_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33128190;  1 drivers
v0x5c7c32d4af30_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c331292e0;  1 drivers
v0x5c7c32d4afd0_0 .net "tmp_sum_out", 0 0, L_0x5c7c33128ce0;  1 drivers
S_0x5c7c32d2ca80 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32d2c880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d38570_0 .net "a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d38720_0 .net "b", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d388f0_0 .net "carry", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d38990_0 .net "sum", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
S_0x5c7c32d2cc60 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d2ca80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d2dd50_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d2de20_0 .net "in_b", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d2def0_0 .net "out", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d2e010_0 .net "temp_out", 0 0, L_0x5c7c32d2b740;  1 drivers
S_0x5c7c32d2ced0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d2cc60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d2b740 .functor NAND 1, L_0x5c7c33125b30, L_0x5c7c3312a560, C4<1>, C4<1>;
v0x5c7c32d2d140_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d2d220_0 .net "in_b", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d2d2e0_0 .net "out", 0 0, L_0x5c7c32d2b740;  alias, 1 drivers
S_0x5c7c32d2d430 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d2cc60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d2dba0_0 .net "in_a", 0 0, L_0x5c7c32d2b740;  alias, 1 drivers
v0x5c7c32d2dc40_0 .net "out", 0 0, L_0x5c7c33128190;  alias, 1 drivers
S_0x5c7c32d2d650 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d2d430;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128190 .functor NAND 1, L_0x5c7c32d2b740, L_0x5c7c32d2b740, C4<1>, C4<1>;
v0x5c7c32d2d8c0_0 .net "in_a", 0 0, L_0x5c7c32d2b740;  alias, 1 drivers
v0x5c7c32d2d9b0_0 .net "in_b", 0 0, L_0x5c7c32d2b740;  alias, 1 drivers
v0x5c7c32d2daa0_0 .net "out", 0 0, L_0x5c7c33128190;  alias, 1 drivers
S_0x5c7c32d2e0d0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d2ca80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d37e90_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d37f30_0 .net "in_b", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d37ff0_0 .net "out", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d38090_0 .net "temp_a_and_out", 0 0, L_0x5c7c331283a0;  1 drivers
v0x5c7c32d38240_0 .net "temp_a_out", 0 0, L_0x5c7c33128240;  1 drivers
v0x5c7c32d382e0_0 .net "temp_b_and_out", 0 0, L_0x5c7c331285b0;  1 drivers
v0x5c7c32d38490_0 .net "temp_b_out", 0 0, L_0x5c7c33128450;  1 drivers
S_0x5c7c32d2e2b0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d2e0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d2f370_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d2f410_0 .net "in_b", 0 0, L_0x5c7c33128240;  alias, 1 drivers
v0x5c7c32d2f500_0 .net "out", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
v0x5c7c32d2f620_0 .net "temp_out", 0 0, L_0x5c7c331282f0;  1 drivers
S_0x5c7c32d2e520 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d2e2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331282f0 .functor NAND 1, L_0x5c7c33125b30, L_0x5c7c33128240, C4<1>, C4<1>;
v0x5c7c32d2e790_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d2e8a0_0 .net "in_b", 0 0, L_0x5c7c33128240;  alias, 1 drivers
v0x5c7c32d2e960_0 .net "out", 0 0, L_0x5c7c331282f0;  alias, 1 drivers
S_0x5c7c32d2ea80 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d2e2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d2f1c0_0 .net "in_a", 0 0, L_0x5c7c331282f0;  alias, 1 drivers
v0x5c7c32d2f260_0 .net "out", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
S_0x5c7c32d2eca0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d2ea80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331283a0 .functor NAND 1, L_0x5c7c331282f0, L_0x5c7c331282f0, C4<1>, C4<1>;
v0x5c7c32d2ef10_0 .net "in_a", 0 0, L_0x5c7c331282f0;  alias, 1 drivers
v0x5c7c32d2efd0_0 .net "in_b", 0 0, L_0x5c7c331282f0;  alias, 1 drivers
v0x5c7c32d2f0c0_0 .net "out", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
S_0x5c7c32d2f6e0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d2e0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d30710_0 .net "in_a", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d307b0_0 .net "in_b", 0 0, L_0x5c7c33128450;  alias, 1 drivers
v0x5c7c32d308a0_0 .net "out", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
v0x5c7c32d309c0_0 .net "temp_out", 0 0, L_0x5c7c33128500;  1 drivers
S_0x5c7c32d2f8c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d2f6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128500 .functor NAND 1, L_0x5c7c3312a560, L_0x5c7c33128450, C4<1>, C4<1>;
v0x5c7c32d2fb30_0 .net "in_a", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d2fc40_0 .net "in_b", 0 0, L_0x5c7c33128450;  alias, 1 drivers
v0x5c7c32d2fd00_0 .net "out", 0 0, L_0x5c7c33128500;  alias, 1 drivers
S_0x5c7c32d2fe20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d2f6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d30560_0 .net "in_a", 0 0, L_0x5c7c33128500;  alias, 1 drivers
v0x5c7c32d30600_0 .net "out", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
S_0x5c7c32d30040 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d2fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331285b0 .functor NAND 1, L_0x5c7c33128500, L_0x5c7c33128500, C4<1>, C4<1>;
v0x5c7c32d302b0_0 .net "in_a", 0 0, L_0x5c7c33128500;  alias, 1 drivers
v0x5c7c32d30370_0 .net "in_b", 0 0, L_0x5c7c33128500;  alias, 1 drivers
v0x5c7c32d30460_0 .net "out", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
S_0x5c7c32d30b10 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d2e0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d31250_0 .net "in_a", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d312f0_0 .net "out", 0 0, L_0x5c7c33128240;  alias, 1 drivers
S_0x5c7c32d30ce0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d30b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128240 .functor NAND 1, L_0x5c7c3312a560, L_0x5c7c3312a560, C4<1>, C4<1>;
v0x5c7c32d30f30_0 .net "in_a", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d31080_0 .net "in_b", 0 0, L_0x5c7c3312a560;  alias, 1 drivers
v0x5c7c32d31140_0 .net "out", 0 0, L_0x5c7c33128240;  alias, 1 drivers
S_0x5c7c32d313f0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d2e0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d31b70_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d31c10_0 .net "out", 0 0, L_0x5c7c33128450;  alias, 1 drivers
S_0x5c7c32d31610 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d313f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128450 .functor NAND 1, L_0x5c7c33125b30, L_0x5c7c33125b30, C4<1>, C4<1>;
v0x5c7c32d31880_0 .net "in_a", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d319d0_0 .net "in_b", 0 0, L_0x5c7c33125b30;  alias, 1 drivers
v0x5c7c32d31a90_0 .net "out", 0 0, L_0x5c7c33128450;  alias, 1 drivers
S_0x5c7c32d31d10 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d2e0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d377e0_0 .net "branch1_out", 0 0, L_0x5c7c331287c0;  1 drivers
v0x5c7c32d37910_0 .net "branch2_out", 0 0, L_0x5c7c33128a50;  1 drivers
v0x5c7c32d37a60_0 .net "in_a", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
v0x5c7c32d37b30_0 .net "in_b", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
v0x5c7c32d37bd0_0 .net "out", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d37c70_0 .net "temp1_out", 0 0, L_0x5c7c33128710;  1 drivers
v0x5c7c32d37d10_0 .net "temp2_out", 0 0, L_0x5c7c331289a0;  1 drivers
v0x5c7c32d37db0_0 .net "temp3_out", 0 0, L_0x5c7c33128c30;  1 drivers
S_0x5c7c32d31f90 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d31d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d33020_0 .net "in_a", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
v0x5c7c32d330c0_0 .net "in_b", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
v0x5c7c32d33180_0 .net "out", 0 0, L_0x5c7c33128710;  alias, 1 drivers
v0x5c7c32d332a0_0 .net "temp_out", 0 0, L_0x5c7c33128660;  1 drivers
S_0x5c7c32d32200 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d31f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128660 .functor NAND 1, L_0x5c7c331283a0, L_0x5c7c331283a0, C4<1>, C4<1>;
v0x5c7c32d32470_0 .net "in_a", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
v0x5c7c32d32530_0 .net "in_b", 0 0, L_0x5c7c331283a0;  alias, 1 drivers
v0x5c7c32d32680_0 .net "out", 0 0, L_0x5c7c33128660;  alias, 1 drivers
S_0x5c7c32d32780 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d31f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d32e70_0 .net "in_a", 0 0, L_0x5c7c33128660;  alias, 1 drivers
v0x5c7c32d32f10_0 .net "out", 0 0, L_0x5c7c33128710;  alias, 1 drivers
S_0x5c7c32d32950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d32780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128710 .functor NAND 1, L_0x5c7c33128660, L_0x5c7c33128660, C4<1>, C4<1>;
v0x5c7c32d32bc0_0 .net "in_a", 0 0, L_0x5c7c33128660;  alias, 1 drivers
v0x5c7c32d32c80_0 .net "in_b", 0 0, L_0x5c7c33128660;  alias, 1 drivers
v0x5c7c32d32d70_0 .net "out", 0 0, L_0x5c7c33128710;  alias, 1 drivers
S_0x5c7c32d33410 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d31d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d34440_0 .net "in_a", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
v0x5c7c32d344e0_0 .net "in_b", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
v0x5c7c32d345a0_0 .net "out", 0 0, L_0x5c7c331289a0;  alias, 1 drivers
v0x5c7c32d346c0_0 .net "temp_out", 0 0, L_0x5c7c32d36260;  1 drivers
S_0x5c7c32d335f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d33410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d36260 .functor NAND 1, L_0x5c7c331285b0, L_0x5c7c331285b0, C4<1>, C4<1>;
v0x5c7c32d33860_0 .net "in_a", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
v0x5c7c32d33920_0 .net "in_b", 0 0, L_0x5c7c331285b0;  alias, 1 drivers
v0x5c7c32d33a70_0 .net "out", 0 0, L_0x5c7c32d36260;  alias, 1 drivers
S_0x5c7c32d33b70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d33410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d34290_0 .net "in_a", 0 0, L_0x5c7c32d36260;  alias, 1 drivers
v0x5c7c32d34330_0 .net "out", 0 0, L_0x5c7c331289a0;  alias, 1 drivers
S_0x5c7c32d33d40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d33b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331289a0 .functor NAND 1, L_0x5c7c32d36260, L_0x5c7c32d36260, C4<1>, C4<1>;
v0x5c7c32d33fb0_0 .net "in_a", 0 0, L_0x5c7c32d36260;  alias, 1 drivers
v0x5c7c32d340a0_0 .net "in_b", 0 0, L_0x5c7c32d36260;  alias, 1 drivers
v0x5c7c32d34190_0 .net "out", 0 0, L_0x5c7c331289a0;  alias, 1 drivers
S_0x5c7c32d34830 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d31d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d35870_0 .net "in_a", 0 0, L_0x5c7c331287c0;  alias, 1 drivers
v0x5c7c32d35940_0 .net "in_b", 0 0, L_0x5c7c33128a50;  alias, 1 drivers
v0x5c7c32d35a10_0 .net "out", 0 0, L_0x5c7c33128c30;  alias, 1 drivers
v0x5c7c32d35b30_0 .net "temp_out", 0 0, L_0x5c7c32d36bd0;  1 drivers
S_0x5c7c32d34a10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d34830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d36bd0 .functor NAND 1, L_0x5c7c331287c0, L_0x5c7c33128a50, C4<1>, C4<1>;
v0x5c7c32d34c60_0 .net "in_a", 0 0, L_0x5c7c331287c0;  alias, 1 drivers
v0x5c7c32d34d40_0 .net "in_b", 0 0, L_0x5c7c33128a50;  alias, 1 drivers
v0x5c7c32d34e00_0 .net "out", 0 0, L_0x5c7c32d36bd0;  alias, 1 drivers
S_0x5c7c32d34f50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d34830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d356c0_0 .net "in_a", 0 0, L_0x5c7c32d36bd0;  alias, 1 drivers
v0x5c7c32d35760_0 .net "out", 0 0, L_0x5c7c33128c30;  alias, 1 drivers
S_0x5c7c32d35170 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d34f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128c30 .functor NAND 1, L_0x5c7c32d36bd0, L_0x5c7c32d36bd0, C4<1>, C4<1>;
v0x5c7c32d353e0_0 .net "in_a", 0 0, L_0x5c7c32d36bd0;  alias, 1 drivers
v0x5c7c32d354d0_0 .net "in_b", 0 0, L_0x5c7c32d36bd0;  alias, 1 drivers
v0x5c7c32d355c0_0 .net "out", 0 0, L_0x5c7c33128c30;  alias, 1 drivers
S_0x5c7c32d35c80 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d31d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d363b0_0 .net "in_a", 0 0, L_0x5c7c33128710;  alias, 1 drivers
v0x5c7c32d36450_0 .net "out", 0 0, L_0x5c7c331287c0;  alias, 1 drivers
S_0x5c7c32d35e50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d35c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331287c0 .functor NAND 1, L_0x5c7c33128710, L_0x5c7c33128710, C4<1>, C4<1>;
v0x5c7c32d360c0_0 .net "in_a", 0 0, L_0x5c7c33128710;  alias, 1 drivers
v0x5c7c32d36180_0 .net "in_b", 0 0, L_0x5c7c33128710;  alias, 1 drivers
v0x5c7c32d362d0_0 .net "out", 0 0, L_0x5c7c331287c0;  alias, 1 drivers
S_0x5c7c32d36550 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d31d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d36d20_0 .net "in_a", 0 0, L_0x5c7c331289a0;  alias, 1 drivers
v0x5c7c32d36dc0_0 .net "out", 0 0, L_0x5c7c33128a50;  alias, 1 drivers
S_0x5c7c32d367c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d36550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128a50 .functor NAND 1, L_0x5c7c331289a0, L_0x5c7c331289a0, C4<1>, C4<1>;
v0x5c7c32d36a30_0 .net "in_a", 0 0, L_0x5c7c331289a0;  alias, 1 drivers
v0x5c7c32d36af0_0 .net "in_b", 0 0, L_0x5c7c331289a0;  alias, 1 drivers
v0x5c7c32d36c40_0 .net "out", 0 0, L_0x5c7c33128a50;  alias, 1 drivers
S_0x5c7c32d36ec0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d31d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d37660_0 .net "in_a", 0 0, L_0x5c7c33128c30;  alias, 1 drivers
v0x5c7c32d37700_0 .net "out", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
S_0x5c7c32d370e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d36ec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33128ce0 .functor NAND 1, L_0x5c7c33128c30, L_0x5c7c33128c30, C4<1>, C4<1>;
v0x5c7c32d37350_0 .net "in_a", 0 0, L_0x5c7c33128c30;  alias, 1 drivers
v0x5c7c32d37410_0 .net "in_b", 0 0, L_0x5c7c33128c30;  alias, 1 drivers
v0x5c7c32d37560_0 .net "out", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
S_0x5c7c32d38a70 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32d2c880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d44520_0 .net "a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d445c0_0 .net "b", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d44680_0 .net "carry", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d44720_0 .net "sum", 0 0, L_0x5c7c33129c10;  alias, 1 drivers
S_0x5c7c32d38c20 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d38a70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d39bc0_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d39c60_0 .net "in_b", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d39d20_0 .net "out", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d39e40_0 .net "temp_out", 0 0, L_0x5c7c32d374f0;  1 drivers
S_0x5c7c32d38dd0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d38c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d374f0 .functor NAND 1, L_0x5c7c33128ce0, L_0x5c7c33127dc0, C4<1>, C4<1>;
v0x5c7c32d39040_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d39100_0 .net "in_b", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d391c0_0 .net "out", 0 0, L_0x5c7c32d374f0;  alias, 1 drivers
S_0x5c7c32d392f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d38c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d39a10_0 .net "in_a", 0 0, L_0x5c7c32d374f0;  alias, 1 drivers
v0x5c7c32d39ab0_0 .net "out", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
S_0x5c7c32d394c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d392f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331292e0 .functor NAND 1, L_0x5c7c32d374f0, L_0x5c7c32d374f0, C4<1>, C4<1>;
v0x5c7c32d39730_0 .net "in_a", 0 0, L_0x5c7c32d374f0;  alias, 1 drivers
v0x5c7c32d39820_0 .net "in_b", 0 0, L_0x5c7c32d374f0;  alias, 1 drivers
v0x5c7c32d39910_0 .net "out", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
S_0x5c7c32d39fb0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d38a70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d43e40_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d43ee0_0 .net "in_b", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d43fa0_0 .net "out", 0 0, L_0x5c7c33129c10;  alias, 1 drivers
v0x5c7c32d44040_0 .net "temp_a_and_out", 0 0, L_0x5c7c331294f0;  1 drivers
v0x5c7c32d441f0_0 .net "temp_a_out", 0 0, L_0x5c7c33129390;  1 drivers
v0x5c7c32d44290_0 .net "temp_b_and_out", 0 0, L_0x5c7c33129700;  1 drivers
v0x5c7c32d44440_0 .net "temp_b_out", 0 0, L_0x5c7c331295a0;  1 drivers
S_0x5c7c32d3a190 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d39fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d3b230_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d3b3e0_0 .net "in_b", 0 0, L_0x5c7c33129390;  alias, 1 drivers
v0x5c7c32d3b4d0_0 .net "out", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
v0x5c7c32d3b5f0_0 .net "temp_out", 0 0, L_0x5c7c33129440;  1 drivers
S_0x5c7c32d3a400 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d3a190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129440 .functor NAND 1, L_0x5c7c33128ce0, L_0x5c7c33129390, C4<1>, C4<1>;
v0x5c7c32d3a670_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d3a730_0 .net "in_b", 0 0, L_0x5c7c33129390;  alias, 1 drivers
v0x5c7c32d3a7f0_0 .net "out", 0 0, L_0x5c7c33129440;  alias, 1 drivers
S_0x5c7c32d3a910 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d3a190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d3b080_0 .net "in_a", 0 0, L_0x5c7c33129440;  alias, 1 drivers
v0x5c7c32d3b120_0 .net "out", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
S_0x5c7c32d3ab30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d3a910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331294f0 .functor NAND 1, L_0x5c7c33129440, L_0x5c7c33129440, C4<1>, C4<1>;
v0x5c7c32d3ada0_0 .net "in_a", 0 0, L_0x5c7c33129440;  alias, 1 drivers
v0x5c7c32d3ae90_0 .net "in_b", 0 0, L_0x5c7c33129440;  alias, 1 drivers
v0x5c7c32d3af80_0 .net "out", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
S_0x5c7c32d3b6b0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d39fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d3c6c0_0 .net "in_a", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d3c760_0 .net "in_b", 0 0, L_0x5c7c331295a0;  alias, 1 drivers
v0x5c7c32d3c850_0 .net "out", 0 0, L_0x5c7c33129700;  alias, 1 drivers
v0x5c7c32d3c970_0 .net "temp_out", 0 0, L_0x5c7c33129650;  1 drivers
S_0x5c7c32d3b890 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d3b6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129650 .functor NAND 1, L_0x5c7c33127dc0, L_0x5c7c331295a0, C4<1>, C4<1>;
v0x5c7c32d3bb00_0 .net "in_a", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d3bbc0_0 .net "in_b", 0 0, L_0x5c7c331295a0;  alias, 1 drivers
v0x5c7c32d3bc80_0 .net "out", 0 0, L_0x5c7c33129650;  alias, 1 drivers
S_0x5c7c32d3bda0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d3b6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d3c510_0 .net "in_a", 0 0, L_0x5c7c33129650;  alias, 1 drivers
v0x5c7c32d3c5b0_0 .net "out", 0 0, L_0x5c7c33129700;  alias, 1 drivers
S_0x5c7c32d3bfc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d3bda0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129700 .functor NAND 1, L_0x5c7c33129650, L_0x5c7c33129650, C4<1>, C4<1>;
v0x5c7c32d3c230_0 .net "in_a", 0 0, L_0x5c7c33129650;  alias, 1 drivers
v0x5c7c32d3c320_0 .net "in_b", 0 0, L_0x5c7c33129650;  alias, 1 drivers
v0x5c7c32d3c410_0 .net "out", 0 0, L_0x5c7c33129700;  alias, 1 drivers
S_0x5c7c32d3cac0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d39fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d3d2d0_0 .net "in_a", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d3d370_0 .net "out", 0 0, L_0x5c7c33129390;  alias, 1 drivers
S_0x5c7c32d3cc90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d3cac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129390 .functor NAND 1, L_0x5c7c33127dc0, L_0x5c7c33127dc0, C4<1>, C4<1>;
v0x5c7c32d3cee0_0 .net "in_a", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d3d0b0_0 .net "in_b", 0 0, L_0x5c7c33127dc0;  alias, 1 drivers
v0x5c7c32d3d170_0 .net "out", 0 0, L_0x5c7c33129390;  alias, 1 drivers
S_0x5c7c32d3d470 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d39fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d3dbb0_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d3dc50_0 .net "out", 0 0, L_0x5c7c331295a0;  alias, 1 drivers
S_0x5c7c32d3d690 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d3d470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331295a0 .functor NAND 1, L_0x5c7c33128ce0, L_0x5c7c33128ce0, C4<1>, C4<1>;
v0x5c7c32d3d900_0 .net "in_a", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d3d9c0_0 .net "in_b", 0 0, L_0x5c7c33128ce0;  alias, 1 drivers
v0x5c7c32d3da80_0 .net "out", 0 0, L_0x5c7c331295a0;  alias, 1 drivers
S_0x5c7c32d3dd50 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d39fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d43790_0 .net "branch1_out", 0 0, L_0x5c7c33129910;  1 drivers
v0x5c7c32d438c0_0 .net "branch2_out", 0 0, L_0x5c7c33129a90;  1 drivers
v0x5c7c32d43a10_0 .net "in_a", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
v0x5c7c32d43ae0_0 .net "in_b", 0 0, L_0x5c7c33129700;  alias, 1 drivers
v0x5c7c32d43b80_0 .net "out", 0 0, L_0x5c7c33129c10;  alias, 1 drivers
v0x5c7c32d43c20_0 .net "temp1_out", 0 0, L_0x5c7c33129860;  1 drivers
v0x5c7c32d43cc0_0 .net "temp2_out", 0 0, L_0x5c7c331299e0;  1 drivers
v0x5c7c32d43d60_0 .net "temp3_out", 0 0, L_0x5c7c33129b60;  1 drivers
S_0x5c7c32d3dfd0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d3dd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d3efd0_0 .net "in_a", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
v0x5c7c32d3f070_0 .net "in_b", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
v0x5c7c32d3f130_0 .net "out", 0 0, L_0x5c7c33129860;  alias, 1 drivers
v0x5c7c32d3f250_0 .net "temp_out", 0 0, L_0x5c7c331297b0;  1 drivers
S_0x5c7c32d3e240 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d3dfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331297b0 .functor NAND 1, L_0x5c7c331294f0, L_0x5c7c331294f0, C4<1>, C4<1>;
v0x5c7c32d3e4b0_0 .net "in_a", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
v0x5c7c32d3e570_0 .net "in_b", 0 0, L_0x5c7c331294f0;  alias, 1 drivers
v0x5c7c32d3e630_0 .net "out", 0 0, L_0x5c7c331297b0;  alias, 1 drivers
S_0x5c7c32d3e730 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d3dfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d3ee20_0 .net "in_a", 0 0, L_0x5c7c331297b0;  alias, 1 drivers
v0x5c7c32d3eec0_0 .net "out", 0 0, L_0x5c7c33129860;  alias, 1 drivers
S_0x5c7c32d3e900 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d3e730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129860 .functor NAND 1, L_0x5c7c331297b0, L_0x5c7c331297b0, C4<1>, C4<1>;
v0x5c7c32d3eb70_0 .net "in_a", 0 0, L_0x5c7c331297b0;  alias, 1 drivers
v0x5c7c32d3ec30_0 .net "in_b", 0 0, L_0x5c7c331297b0;  alias, 1 drivers
v0x5c7c32d3ed20_0 .net "out", 0 0, L_0x5c7c33129860;  alias, 1 drivers
S_0x5c7c32d3f3c0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d3dd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d403f0_0 .net "in_a", 0 0, L_0x5c7c33129700;  alias, 1 drivers
v0x5c7c32d40490_0 .net "in_b", 0 0, L_0x5c7c33129700;  alias, 1 drivers
v0x5c7c32d40550_0 .net "out", 0 0, L_0x5c7c331299e0;  alias, 1 drivers
v0x5c7c32d40670_0 .net "temp_out", 0 0, L_0x5c7c32d42210;  1 drivers
S_0x5c7c32d3f5a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d3f3c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d42210 .functor NAND 1, L_0x5c7c33129700, L_0x5c7c33129700, C4<1>, C4<1>;
v0x5c7c32d3f810_0 .net "in_a", 0 0, L_0x5c7c33129700;  alias, 1 drivers
v0x5c7c32d3f8d0_0 .net "in_b", 0 0, L_0x5c7c33129700;  alias, 1 drivers
v0x5c7c32d3fa20_0 .net "out", 0 0, L_0x5c7c32d42210;  alias, 1 drivers
S_0x5c7c32d3fb20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d3f3c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d40240_0 .net "in_a", 0 0, L_0x5c7c32d42210;  alias, 1 drivers
v0x5c7c32d402e0_0 .net "out", 0 0, L_0x5c7c331299e0;  alias, 1 drivers
S_0x5c7c32d3fcf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d3fb20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331299e0 .functor NAND 1, L_0x5c7c32d42210, L_0x5c7c32d42210, C4<1>, C4<1>;
v0x5c7c32d3ff60_0 .net "in_a", 0 0, L_0x5c7c32d42210;  alias, 1 drivers
v0x5c7c32d40050_0 .net "in_b", 0 0, L_0x5c7c32d42210;  alias, 1 drivers
v0x5c7c32d40140_0 .net "out", 0 0, L_0x5c7c331299e0;  alias, 1 drivers
S_0x5c7c32d407e0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d3dd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d41820_0 .net "in_a", 0 0, L_0x5c7c33129910;  alias, 1 drivers
v0x5c7c32d418f0_0 .net "in_b", 0 0, L_0x5c7c33129a90;  alias, 1 drivers
v0x5c7c32d419c0_0 .net "out", 0 0, L_0x5c7c33129b60;  alias, 1 drivers
v0x5c7c32d41ae0_0 .net "temp_out", 0 0, L_0x5c7c32d42b80;  1 drivers
S_0x5c7c32d409c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d407e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d42b80 .functor NAND 1, L_0x5c7c33129910, L_0x5c7c33129a90, C4<1>, C4<1>;
v0x5c7c32d40c10_0 .net "in_a", 0 0, L_0x5c7c33129910;  alias, 1 drivers
v0x5c7c32d40cf0_0 .net "in_b", 0 0, L_0x5c7c33129a90;  alias, 1 drivers
v0x5c7c32d40db0_0 .net "out", 0 0, L_0x5c7c32d42b80;  alias, 1 drivers
S_0x5c7c32d40f00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d407e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d41670_0 .net "in_a", 0 0, L_0x5c7c32d42b80;  alias, 1 drivers
v0x5c7c32d41710_0 .net "out", 0 0, L_0x5c7c33129b60;  alias, 1 drivers
S_0x5c7c32d41120 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d40f00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129b60 .functor NAND 1, L_0x5c7c32d42b80, L_0x5c7c32d42b80, C4<1>, C4<1>;
v0x5c7c32d41390_0 .net "in_a", 0 0, L_0x5c7c32d42b80;  alias, 1 drivers
v0x5c7c32d41480_0 .net "in_b", 0 0, L_0x5c7c32d42b80;  alias, 1 drivers
v0x5c7c32d41570_0 .net "out", 0 0, L_0x5c7c33129b60;  alias, 1 drivers
S_0x5c7c32d41c30 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d3dd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d42360_0 .net "in_a", 0 0, L_0x5c7c33129860;  alias, 1 drivers
v0x5c7c32d42400_0 .net "out", 0 0, L_0x5c7c33129910;  alias, 1 drivers
S_0x5c7c32d41e00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d41c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129910 .functor NAND 1, L_0x5c7c33129860, L_0x5c7c33129860, C4<1>, C4<1>;
v0x5c7c32d42070_0 .net "in_a", 0 0, L_0x5c7c33129860;  alias, 1 drivers
v0x5c7c32d42130_0 .net "in_b", 0 0, L_0x5c7c33129860;  alias, 1 drivers
v0x5c7c32d42280_0 .net "out", 0 0, L_0x5c7c33129910;  alias, 1 drivers
S_0x5c7c32d42500 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d3dd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d42cd0_0 .net "in_a", 0 0, L_0x5c7c331299e0;  alias, 1 drivers
v0x5c7c32d42d70_0 .net "out", 0 0, L_0x5c7c33129a90;  alias, 1 drivers
S_0x5c7c32d42770 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d42500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129a90 .functor NAND 1, L_0x5c7c331299e0, L_0x5c7c331299e0, C4<1>, C4<1>;
v0x5c7c32d429e0_0 .net "in_a", 0 0, L_0x5c7c331299e0;  alias, 1 drivers
v0x5c7c32d42aa0_0 .net "in_b", 0 0, L_0x5c7c331299e0;  alias, 1 drivers
v0x5c7c32d42bf0_0 .net "out", 0 0, L_0x5c7c33129a90;  alias, 1 drivers
S_0x5c7c32d42e70 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d3dd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d43610_0 .net "in_a", 0 0, L_0x5c7c33129b60;  alias, 1 drivers
v0x5c7c32d436b0_0 .net "out", 0 0, L_0x5c7c33129c10;  alias, 1 drivers
S_0x5c7c32d43090 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d42e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129c10 .functor NAND 1, L_0x5c7c33129b60, L_0x5c7c33129b60, C4<1>, C4<1>;
v0x5c7c32d43300_0 .net "in_a", 0 0, L_0x5c7c33129b60;  alias, 1 drivers
v0x5c7c32d433c0_0 .net "in_b", 0 0, L_0x5c7c33129b60;  alias, 1 drivers
v0x5c7c32d43510_0 .net "out", 0 0, L_0x5c7c33129c10;  alias, 1 drivers
S_0x5c7c32d44890 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32d2c880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d4a280_0 .net "branch1_out", 0 0, L_0x5c7c33129ea0;  1 drivers
v0x5c7c32d4a3b0_0 .net "branch2_out", 0 0, L_0x5c7c3312a130;  1 drivers
v0x5c7c32d4a500_0 .net "in_a", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d4a6e0_0 .net "in_b", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d4a890_0 .net "out", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d4a930_0 .net "temp1_out", 0 0, L_0x5c7c33129df0;  1 drivers
v0x5c7c32d4a9d0_0 .net "temp2_out", 0 0, L_0x5c7c3312a080;  1 drivers
v0x5c7c32d4aa70_0 .net "temp3_out", 0 0, L_0x5c7c3312a310;  1 drivers
S_0x5c7c32d44a20 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d44890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d45ac0_0 .net "in_a", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d45b60_0 .net "in_b", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d45c20_0 .net "out", 0 0, L_0x5c7c33129df0;  alias, 1 drivers
v0x5c7c32d45d40_0 .net "temp_out", 0 0, L_0x5c7c32d434a0;  1 drivers
S_0x5c7c32d44c40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d44a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d434a0 .functor NAND 1, L_0x5c7c33128190, L_0x5c7c33128190, C4<1>, C4<1>;
v0x5c7c32d44eb0_0 .net "in_a", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d45000_0 .net "in_b", 0 0, L_0x5c7c33128190;  alias, 1 drivers
v0x5c7c32d450c0_0 .net "out", 0 0, L_0x5c7c32d434a0;  alias, 1 drivers
S_0x5c7c32d451f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d44a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d45910_0 .net "in_a", 0 0, L_0x5c7c32d434a0;  alias, 1 drivers
v0x5c7c32d459b0_0 .net "out", 0 0, L_0x5c7c33129df0;  alias, 1 drivers
S_0x5c7c32d453c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d451f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129df0 .functor NAND 1, L_0x5c7c32d434a0, L_0x5c7c32d434a0, C4<1>, C4<1>;
v0x5c7c32d45630_0 .net "in_a", 0 0, L_0x5c7c32d434a0;  alias, 1 drivers
v0x5c7c32d45720_0 .net "in_b", 0 0, L_0x5c7c32d434a0;  alias, 1 drivers
v0x5c7c32d45810_0 .net "out", 0 0, L_0x5c7c33129df0;  alias, 1 drivers
S_0x5c7c32d45eb0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d44890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d46ee0_0 .net "in_a", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d46f80_0 .net "in_b", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d47040_0 .net "out", 0 0, L_0x5c7c3312a080;  alias, 1 drivers
v0x5c7c32d47160_0 .net "temp_out", 0 0, L_0x5c7c32d48d00;  1 drivers
S_0x5c7c32d46090 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d45eb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d48d00 .functor NAND 1, L_0x5c7c331292e0, L_0x5c7c331292e0, C4<1>, C4<1>;
v0x5c7c32d46300_0 .net "in_a", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d46450_0 .net "in_b", 0 0, L_0x5c7c331292e0;  alias, 1 drivers
v0x5c7c32d46510_0 .net "out", 0 0, L_0x5c7c32d48d00;  alias, 1 drivers
S_0x5c7c32d46610 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d45eb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d46d30_0 .net "in_a", 0 0, L_0x5c7c32d48d00;  alias, 1 drivers
v0x5c7c32d46dd0_0 .net "out", 0 0, L_0x5c7c3312a080;  alias, 1 drivers
S_0x5c7c32d467e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d46610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a080 .functor NAND 1, L_0x5c7c32d48d00, L_0x5c7c32d48d00, C4<1>, C4<1>;
v0x5c7c32d46a50_0 .net "in_a", 0 0, L_0x5c7c32d48d00;  alias, 1 drivers
v0x5c7c32d46b40_0 .net "in_b", 0 0, L_0x5c7c32d48d00;  alias, 1 drivers
v0x5c7c32d46c30_0 .net "out", 0 0, L_0x5c7c3312a080;  alias, 1 drivers
S_0x5c7c32d472d0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d44890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d48310_0 .net "in_a", 0 0, L_0x5c7c33129ea0;  alias, 1 drivers
v0x5c7c32d483e0_0 .net "in_b", 0 0, L_0x5c7c3312a130;  alias, 1 drivers
v0x5c7c32d484b0_0 .net "out", 0 0, L_0x5c7c3312a310;  alias, 1 drivers
v0x5c7c32d485d0_0 .net "temp_out", 0 0, L_0x5c7c32d49670;  1 drivers
S_0x5c7c32d474b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d472d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d49670 .functor NAND 1, L_0x5c7c33129ea0, L_0x5c7c3312a130, C4<1>, C4<1>;
v0x5c7c32d47700_0 .net "in_a", 0 0, L_0x5c7c33129ea0;  alias, 1 drivers
v0x5c7c32d477e0_0 .net "in_b", 0 0, L_0x5c7c3312a130;  alias, 1 drivers
v0x5c7c32d478a0_0 .net "out", 0 0, L_0x5c7c32d49670;  alias, 1 drivers
S_0x5c7c32d479f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d472d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d48160_0 .net "in_a", 0 0, L_0x5c7c32d49670;  alias, 1 drivers
v0x5c7c32d48200_0 .net "out", 0 0, L_0x5c7c3312a310;  alias, 1 drivers
S_0x5c7c32d47c10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d479f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a310 .functor NAND 1, L_0x5c7c32d49670, L_0x5c7c32d49670, C4<1>, C4<1>;
v0x5c7c32d47e80_0 .net "in_a", 0 0, L_0x5c7c32d49670;  alias, 1 drivers
v0x5c7c32d47f70_0 .net "in_b", 0 0, L_0x5c7c32d49670;  alias, 1 drivers
v0x5c7c32d48060_0 .net "out", 0 0, L_0x5c7c3312a310;  alias, 1 drivers
S_0x5c7c32d48720 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d44890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d48e50_0 .net "in_a", 0 0, L_0x5c7c33129df0;  alias, 1 drivers
v0x5c7c32d48ef0_0 .net "out", 0 0, L_0x5c7c33129ea0;  alias, 1 drivers
S_0x5c7c32d488f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d48720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33129ea0 .functor NAND 1, L_0x5c7c33129df0, L_0x5c7c33129df0, C4<1>, C4<1>;
v0x5c7c32d48b60_0 .net "in_a", 0 0, L_0x5c7c33129df0;  alias, 1 drivers
v0x5c7c32d48c20_0 .net "in_b", 0 0, L_0x5c7c33129df0;  alias, 1 drivers
v0x5c7c32d48d70_0 .net "out", 0 0, L_0x5c7c33129ea0;  alias, 1 drivers
S_0x5c7c32d48ff0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d44890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d497c0_0 .net "in_a", 0 0, L_0x5c7c3312a080;  alias, 1 drivers
v0x5c7c32d49860_0 .net "out", 0 0, L_0x5c7c3312a130;  alias, 1 drivers
S_0x5c7c32d49260 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d48ff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a130 .functor NAND 1, L_0x5c7c3312a080, L_0x5c7c3312a080, C4<1>, C4<1>;
v0x5c7c32d494d0_0 .net "in_a", 0 0, L_0x5c7c3312a080;  alias, 1 drivers
v0x5c7c32d49590_0 .net "in_b", 0 0, L_0x5c7c3312a080;  alias, 1 drivers
v0x5c7c32d496e0_0 .net "out", 0 0, L_0x5c7c3312a130;  alias, 1 drivers
S_0x5c7c32d49960 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d44890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d4a100_0 .net "in_a", 0 0, L_0x5c7c3312a310;  alias, 1 drivers
v0x5c7c32d4a1a0_0 .net "out", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
S_0x5c7c32d49b80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d49960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a3c0 .functor NAND 1, L_0x5c7c3312a310, L_0x5c7c3312a310, C4<1>, C4<1>;
v0x5c7c32d49df0_0 .net "in_a", 0 0, L_0x5c7c3312a310;  alias, 1 drivers
v0x5c7c32d49eb0_0 .net "in_b", 0 0, L_0x5c7c3312a310;  alias, 1 drivers
v0x5c7c32d4a000_0 .net "out", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
S_0x5c7c32d4b0d0 .scope module, "fa_gate12" "FullAdder" 2 17, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32d693b0_0 .net "a", 0 0, L_0x5c7c3312cad0;  1 drivers
v0x5c7c32d69450_0 .net "b", 0 0, L_0x5c7c3312cb70;  1 drivers
v0x5c7c32d69510_0 .net "c", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d695b0_0 .net "carry", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d69650_0 .net "sum", 0 0, L_0x5c7c3312c180;  1 drivers
v0x5c7c32d696f0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c3312a700;  1 drivers
v0x5c7c32d69790_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c3312b850;  1 drivers
v0x5c7c32d69830_0 .net "tmp_sum_out", 0 0, L_0x5c7c3312b250;  1 drivers
S_0x5c7c32d4b2b0 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32d4b0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d56dd0_0 .net "a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d56f80_0 .net "b", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d57150_0 .net "carry", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d571f0_0 .net "sum", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
S_0x5c7c32d4b4c0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d4b2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d4c5b0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d4c680_0 .net "in_b", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4c750_0 .net "out", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d4c870_0 .net "temp_out", 0 0, L_0x5c7c32d49f90;  1 drivers
S_0x5c7c32d4b730 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d4b4c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d49f90 .functor NAND 1, L_0x5c7c3312cad0, L_0x5c7c3312cb70, C4<1>, C4<1>;
v0x5c7c32d4b9a0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d4ba80_0 .net "in_b", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4bb40_0 .net "out", 0 0, L_0x5c7c32d49f90;  alias, 1 drivers
S_0x5c7c32d4bc90 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d4b4c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d4c400_0 .net "in_a", 0 0, L_0x5c7c32d49f90;  alias, 1 drivers
v0x5c7c32d4c4a0_0 .net "out", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
S_0x5c7c32d4beb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d4bc90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a700 .functor NAND 1, L_0x5c7c32d49f90, L_0x5c7c32d49f90, C4<1>, C4<1>;
v0x5c7c32d4c120_0 .net "in_a", 0 0, L_0x5c7c32d49f90;  alias, 1 drivers
v0x5c7c32d4c210_0 .net "in_b", 0 0, L_0x5c7c32d49f90;  alias, 1 drivers
v0x5c7c32d4c300_0 .net "out", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
S_0x5c7c32d4c930 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d4b2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d566f0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d56790_0 .net "in_b", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d56850_0 .net "out", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d568f0_0 .net "temp_a_and_out", 0 0, L_0x5c7c3312a910;  1 drivers
v0x5c7c32d56aa0_0 .net "temp_a_out", 0 0, L_0x5c7c3312a7b0;  1 drivers
v0x5c7c32d56b40_0 .net "temp_b_and_out", 0 0, L_0x5c7c3312ab20;  1 drivers
v0x5c7c32d56cf0_0 .net "temp_b_out", 0 0, L_0x5c7c3312a9c0;  1 drivers
S_0x5c7c32d4cb10 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d4c930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d4dbd0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d4dc70_0 .net "in_b", 0 0, L_0x5c7c3312a7b0;  alias, 1 drivers
v0x5c7c32d4dd60_0 .net "out", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
v0x5c7c32d4de80_0 .net "temp_out", 0 0, L_0x5c7c3312a860;  1 drivers
S_0x5c7c32d4cd80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d4cb10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a860 .functor NAND 1, L_0x5c7c3312cad0, L_0x5c7c3312a7b0, C4<1>, C4<1>;
v0x5c7c32d4cff0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d4d100_0 .net "in_b", 0 0, L_0x5c7c3312a7b0;  alias, 1 drivers
v0x5c7c32d4d1c0_0 .net "out", 0 0, L_0x5c7c3312a860;  alias, 1 drivers
S_0x5c7c32d4d2e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d4cb10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d4da20_0 .net "in_a", 0 0, L_0x5c7c3312a860;  alias, 1 drivers
v0x5c7c32d4dac0_0 .net "out", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
S_0x5c7c32d4d500 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d4d2e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a910 .functor NAND 1, L_0x5c7c3312a860, L_0x5c7c3312a860, C4<1>, C4<1>;
v0x5c7c32d4d770_0 .net "in_a", 0 0, L_0x5c7c3312a860;  alias, 1 drivers
v0x5c7c32d4d830_0 .net "in_b", 0 0, L_0x5c7c3312a860;  alias, 1 drivers
v0x5c7c32d4d920_0 .net "out", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
S_0x5c7c32d4df40 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d4c930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d4ef70_0 .net "in_a", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4f010_0 .net "in_b", 0 0, L_0x5c7c3312a9c0;  alias, 1 drivers
v0x5c7c32d4f100_0 .net "out", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
v0x5c7c32d4f220_0 .net "temp_out", 0 0, L_0x5c7c3312aa70;  1 drivers
S_0x5c7c32d4e120 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d4df40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312aa70 .functor NAND 1, L_0x5c7c3312cb70, L_0x5c7c3312a9c0, C4<1>, C4<1>;
v0x5c7c32d4e390_0 .net "in_a", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4e4a0_0 .net "in_b", 0 0, L_0x5c7c3312a9c0;  alias, 1 drivers
v0x5c7c32d4e560_0 .net "out", 0 0, L_0x5c7c3312aa70;  alias, 1 drivers
S_0x5c7c32d4e680 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d4df40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d4edc0_0 .net "in_a", 0 0, L_0x5c7c3312aa70;  alias, 1 drivers
v0x5c7c32d4ee60_0 .net "out", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
S_0x5c7c32d4e8a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d4e680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ab20 .functor NAND 1, L_0x5c7c3312aa70, L_0x5c7c3312aa70, C4<1>, C4<1>;
v0x5c7c32d4eb10_0 .net "in_a", 0 0, L_0x5c7c3312aa70;  alias, 1 drivers
v0x5c7c32d4ebd0_0 .net "in_b", 0 0, L_0x5c7c3312aa70;  alias, 1 drivers
v0x5c7c32d4ecc0_0 .net "out", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
S_0x5c7c32d4f370 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d4c930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d4fab0_0 .net "in_a", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4fb50_0 .net "out", 0 0, L_0x5c7c3312a7b0;  alias, 1 drivers
S_0x5c7c32d4f540 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d4f370;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a7b0 .functor NAND 1, L_0x5c7c3312cb70, L_0x5c7c3312cb70, C4<1>, C4<1>;
v0x5c7c32d4f790_0 .net "in_a", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4f8e0_0 .net "in_b", 0 0, L_0x5c7c3312cb70;  alias, 1 drivers
v0x5c7c32d4f9a0_0 .net "out", 0 0, L_0x5c7c3312a7b0;  alias, 1 drivers
S_0x5c7c32d4fc50 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d4c930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d503d0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d50470_0 .net "out", 0 0, L_0x5c7c3312a9c0;  alias, 1 drivers
S_0x5c7c32d4fe70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d4fc50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312a9c0 .functor NAND 1, L_0x5c7c3312cad0, L_0x5c7c3312cad0, C4<1>, C4<1>;
v0x5c7c32d500e0_0 .net "in_a", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d50230_0 .net "in_b", 0 0, L_0x5c7c3312cad0;  alias, 1 drivers
v0x5c7c32d502f0_0 .net "out", 0 0, L_0x5c7c3312a9c0;  alias, 1 drivers
S_0x5c7c32d50570 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d4c930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d56040_0 .net "branch1_out", 0 0, L_0x5c7c3312ad30;  1 drivers
v0x5c7c32d56170_0 .net "branch2_out", 0 0, L_0x5c7c3312afc0;  1 drivers
v0x5c7c32d562c0_0 .net "in_a", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
v0x5c7c32d56390_0 .net "in_b", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
v0x5c7c32d56430_0 .net "out", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d564d0_0 .net "temp1_out", 0 0, L_0x5c7c3312ac80;  1 drivers
v0x5c7c32d56570_0 .net "temp2_out", 0 0, L_0x5c7c3312af10;  1 drivers
v0x5c7c32d56610_0 .net "temp3_out", 0 0, L_0x5c7c3312b1a0;  1 drivers
S_0x5c7c32d507f0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d50570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d51880_0 .net "in_a", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
v0x5c7c32d51920_0 .net "in_b", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
v0x5c7c32d519e0_0 .net "out", 0 0, L_0x5c7c3312ac80;  alias, 1 drivers
v0x5c7c32d51b00_0 .net "temp_out", 0 0, L_0x5c7c3312abd0;  1 drivers
S_0x5c7c32d50a60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d507f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312abd0 .functor NAND 1, L_0x5c7c3312a910, L_0x5c7c3312a910, C4<1>, C4<1>;
v0x5c7c32d50cd0_0 .net "in_a", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
v0x5c7c32d50d90_0 .net "in_b", 0 0, L_0x5c7c3312a910;  alias, 1 drivers
v0x5c7c32d50ee0_0 .net "out", 0 0, L_0x5c7c3312abd0;  alias, 1 drivers
S_0x5c7c32d50fe0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d507f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d516d0_0 .net "in_a", 0 0, L_0x5c7c3312abd0;  alias, 1 drivers
v0x5c7c32d51770_0 .net "out", 0 0, L_0x5c7c3312ac80;  alias, 1 drivers
S_0x5c7c32d511b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d50fe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ac80 .functor NAND 1, L_0x5c7c3312abd0, L_0x5c7c3312abd0, C4<1>, C4<1>;
v0x5c7c32d51420_0 .net "in_a", 0 0, L_0x5c7c3312abd0;  alias, 1 drivers
v0x5c7c32d514e0_0 .net "in_b", 0 0, L_0x5c7c3312abd0;  alias, 1 drivers
v0x5c7c32d515d0_0 .net "out", 0 0, L_0x5c7c3312ac80;  alias, 1 drivers
S_0x5c7c32d51c70 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d50570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d52ca0_0 .net "in_a", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
v0x5c7c32d52d40_0 .net "in_b", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
v0x5c7c32d52e00_0 .net "out", 0 0, L_0x5c7c3312af10;  alias, 1 drivers
v0x5c7c32d52f20_0 .net "temp_out", 0 0, L_0x5c7c32d54ac0;  1 drivers
S_0x5c7c32d51e50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d51c70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d54ac0 .functor NAND 1, L_0x5c7c3312ab20, L_0x5c7c3312ab20, C4<1>, C4<1>;
v0x5c7c32d520c0_0 .net "in_a", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
v0x5c7c32d52180_0 .net "in_b", 0 0, L_0x5c7c3312ab20;  alias, 1 drivers
v0x5c7c32d522d0_0 .net "out", 0 0, L_0x5c7c32d54ac0;  alias, 1 drivers
S_0x5c7c32d523d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d51c70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d52af0_0 .net "in_a", 0 0, L_0x5c7c32d54ac0;  alias, 1 drivers
v0x5c7c32d52b90_0 .net "out", 0 0, L_0x5c7c3312af10;  alias, 1 drivers
S_0x5c7c32d525a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d523d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312af10 .functor NAND 1, L_0x5c7c32d54ac0, L_0x5c7c32d54ac0, C4<1>, C4<1>;
v0x5c7c32d52810_0 .net "in_a", 0 0, L_0x5c7c32d54ac0;  alias, 1 drivers
v0x5c7c32d52900_0 .net "in_b", 0 0, L_0x5c7c32d54ac0;  alias, 1 drivers
v0x5c7c32d529f0_0 .net "out", 0 0, L_0x5c7c3312af10;  alias, 1 drivers
S_0x5c7c32d53090 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d50570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d540d0_0 .net "in_a", 0 0, L_0x5c7c3312ad30;  alias, 1 drivers
v0x5c7c32d541a0_0 .net "in_b", 0 0, L_0x5c7c3312afc0;  alias, 1 drivers
v0x5c7c32d54270_0 .net "out", 0 0, L_0x5c7c3312b1a0;  alias, 1 drivers
v0x5c7c32d54390_0 .net "temp_out", 0 0, L_0x5c7c32d55430;  1 drivers
S_0x5c7c32d53270 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d53090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d55430 .functor NAND 1, L_0x5c7c3312ad30, L_0x5c7c3312afc0, C4<1>, C4<1>;
v0x5c7c32d534c0_0 .net "in_a", 0 0, L_0x5c7c3312ad30;  alias, 1 drivers
v0x5c7c32d535a0_0 .net "in_b", 0 0, L_0x5c7c3312afc0;  alias, 1 drivers
v0x5c7c32d53660_0 .net "out", 0 0, L_0x5c7c32d55430;  alias, 1 drivers
S_0x5c7c32d537b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d53090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d53f20_0 .net "in_a", 0 0, L_0x5c7c32d55430;  alias, 1 drivers
v0x5c7c32d53fc0_0 .net "out", 0 0, L_0x5c7c3312b1a0;  alias, 1 drivers
S_0x5c7c32d539d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d537b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312b1a0 .functor NAND 1, L_0x5c7c32d55430, L_0x5c7c32d55430, C4<1>, C4<1>;
v0x5c7c32d53c40_0 .net "in_a", 0 0, L_0x5c7c32d55430;  alias, 1 drivers
v0x5c7c32d53d30_0 .net "in_b", 0 0, L_0x5c7c32d55430;  alias, 1 drivers
v0x5c7c32d53e20_0 .net "out", 0 0, L_0x5c7c3312b1a0;  alias, 1 drivers
S_0x5c7c32d544e0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d50570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d54c10_0 .net "in_a", 0 0, L_0x5c7c3312ac80;  alias, 1 drivers
v0x5c7c32d54cb0_0 .net "out", 0 0, L_0x5c7c3312ad30;  alias, 1 drivers
S_0x5c7c32d546b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d544e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ad30 .functor NAND 1, L_0x5c7c3312ac80, L_0x5c7c3312ac80, C4<1>, C4<1>;
v0x5c7c32d54920_0 .net "in_a", 0 0, L_0x5c7c3312ac80;  alias, 1 drivers
v0x5c7c32d549e0_0 .net "in_b", 0 0, L_0x5c7c3312ac80;  alias, 1 drivers
v0x5c7c32d54b30_0 .net "out", 0 0, L_0x5c7c3312ad30;  alias, 1 drivers
S_0x5c7c32d54db0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d50570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d55580_0 .net "in_a", 0 0, L_0x5c7c3312af10;  alias, 1 drivers
v0x5c7c32d55620_0 .net "out", 0 0, L_0x5c7c3312afc0;  alias, 1 drivers
S_0x5c7c32d55020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d54db0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312afc0 .functor NAND 1, L_0x5c7c3312af10, L_0x5c7c3312af10, C4<1>, C4<1>;
v0x5c7c32d55290_0 .net "in_a", 0 0, L_0x5c7c3312af10;  alias, 1 drivers
v0x5c7c32d55350_0 .net "in_b", 0 0, L_0x5c7c3312af10;  alias, 1 drivers
v0x5c7c32d554a0_0 .net "out", 0 0, L_0x5c7c3312afc0;  alias, 1 drivers
S_0x5c7c32d55720 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d50570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d55ec0_0 .net "in_a", 0 0, L_0x5c7c3312b1a0;  alias, 1 drivers
v0x5c7c32d55f60_0 .net "out", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
S_0x5c7c32d55940 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d55720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312b250 .functor NAND 1, L_0x5c7c3312b1a0, L_0x5c7c3312b1a0, C4<1>, C4<1>;
v0x5c7c32d55bb0_0 .net "in_a", 0 0, L_0x5c7c3312b1a0;  alias, 1 drivers
v0x5c7c32d55c70_0 .net "in_b", 0 0, L_0x5c7c3312b1a0;  alias, 1 drivers
v0x5c7c32d55dc0_0 .net "out", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
S_0x5c7c32d572d0 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32d4b0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d62d80_0 .net "a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d62e20_0 .net "b", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d62ee0_0 .net "carry", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d62f80_0 .net "sum", 0 0, L_0x5c7c3312c180;  alias, 1 drivers
S_0x5c7c32d57480 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d572d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d58420_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d584c0_0 .net "in_b", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d58580_0 .net "out", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d586a0_0 .net "temp_out", 0 0, L_0x5c7c32d55d50;  1 drivers
S_0x5c7c32d57630 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d57480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d55d50 .functor NAND 1, L_0x5c7c3312b250, L_0x5c7c3312a3c0, C4<1>, C4<1>;
v0x5c7c32d578a0_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d57960_0 .net "in_b", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d57a20_0 .net "out", 0 0, L_0x5c7c32d55d50;  alias, 1 drivers
S_0x5c7c32d57b50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d57480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d58270_0 .net "in_a", 0 0, L_0x5c7c32d55d50;  alias, 1 drivers
v0x5c7c32d58310_0 .net "out", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
S_0x5c7c32d57d20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d57b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312b850 .functor NAND 1, L_0x5c7c32d55d50, L_0x5c7c32d55d50, C4<1>, C4<1>;
v0x5c7c32d57f90_0 .net "in_a", 0 0, L_0x5c7c32d55d50;  alias, 1 drivers
v0x5c7c32d58080_0 .net "in_b", 0 0, L_0x5c7c32d55d50;  alias, 1 drivers
v0x5c7c32d58170_0 .net "out", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
S_0x5c7c32d58810 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d572d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d626a0_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d62740_0 .net "in_b", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d62800_0 .net "out", 0 0, L_0x5c7c3312c180;  alias, 1 drivers
v0x5c7c32d628a0_0 .net "temp_a_and_out", 0 0, L_0x5c7c3312ba60;  1 drivers
v0x5c7c32d62a50_0 .net "temp_a_out", 0 0, L_0x5c7c3312b900;  1 drivers
v0x5c7c32d62af0_0 .net "temp_b_and_out", 0 0, L_0x5c7c3312bc70;  1 drivers
v0x5c7c32d62ca0_0 .net "temp_b_out", 0 0, L_0x5c7c3312bb10;  1 drivers
S_0x5c7c32d589f0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d58810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d59a90_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d59c40_0 .net "in_b", 0 0, L_0x5c7c3312b900;  alias, 1 drivers
v0x5c7c32d59d30_0 .net "out", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
v0x5c7c32d59e50_0 .net "temp_out", 0 0, L_0x5c7c3312b9b0;  1 drivers
S_0x5c7c32d58c60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d589f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312b9b0 .functor NAND 1, L_0x5c7c3312b250, L_0x5c7c3312b900, C4<1>, C4<1>;
v0x5c7c32d58ed0_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d58f90_0 .net "in_b", 0 0, L_0x5c7c3312b900;  alias, 1 drivers
v0x5c7c32d59050_0 .net "out", 0 0, L_0x5c7c3312b9b0;  alias, 1 drivers
S_0x5c7c32d59170 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d589f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d598e0_0 .net "in_a", 0 0, L_0x5c7c3312b9b0;  alias, 1 drivers
v0x5c7c32d59980_0 .net "out", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
S_0x5c7c32d59390 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d59170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ba60 .functor NAND 1, L_0x5c7c3312b9b0, L_0x5c7c3312b9b0, C4<1>, C4<1>;
v0x5c7c32d59600_0 .net "in_a", 0 0, L_0x5c7c3312b9b0;  alias, 1 drivers
v0x5c7c32d596f0_0 .net "in_b", 0 0, L_0x5c7c3312b9b0;  alias, 1 drivers
v0x5c7c32d597e0_0 .net "out", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
S_0x5c7c32d59f10 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d58810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d5af20_0 .net "in_a", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d5afc0_0 .net "in_b", 0 0, L_0x5c7c3312bb10;  alias, 1 drivers
v0x5c7c32d5b0b0_0 .net "out", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
v0x5c7c32d5b1d0_0 .net "temp_out", 0 0, L_0x5c7c3312bbc0;  1 drivers
S_0x5c7c32d5a0f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d59f10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312bbc0 .functor NAND 1, L_0x5c7c3312a3c0, L_0x5c7c3312bb10, C4<1>, C4<1>;
v0x5c7c32d5a360_0 .net "in_a", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d5a420_0 .net "in_b", 0 0, L_0x5c7c3312bb10;  alias, 1 drivers
v0x5c7c32d5a4e0_0 .net "out", 0 0, L_0x5c7c3312bbc0;  alias, 1 drivers
S_0x5c7c32d5a600 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d59f10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d5ad70_0 .net "in_a", 0 0, L_0x5c7c3312bbc0;  alias, 1 drivers
v0x5c7c32d5ae10_0 .net "out", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
S_0x5c7c32d5a820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d5a600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312bc70 .functor NAND 1, L_0x5c7c3312bbc0, L_0x5c7c3312bbc0, C4<1>, C4<1>;
v0x5c7c32d5aa90_0 .net "in_a", 0 0, L_0x5c7c3312bbc0;  alias, 1 drivers
v0x5c7c32d5ab80_0 .net "in_b", 0 0, L_0x5c7c3312bbc0;  alias, 1 drivers
v0x5c7c32d5ac70_0 .net "out", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
S_0x5c7c32d5b320 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d58810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d5bb30_0 .net "in_a", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d5bbd0_0 .net "out", 0 0, L_0x5c7c3312b900;  alias, 1 drivers
S_0x5c7c32d5b4f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d5b320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312b900 .functor NAND 1, L_0x5c7c3312a3c0, L_0x5c7c3312a3c0, C4<1>, C4<1>;
v0x5c7c32d5b740_0 .net "in_a", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d5b910_0 .net "in_b", 0 0, L_0x5c7c3312a3c0;  alias, 1 drivers
v0x5c7c32d5b9d0_0 .net "out", 0 0, L_0x5c7c3312b900;  alias, 1 drivers
S_0x5c7c32d5bcd0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d58810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d5c410_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d5c4b0_0 .net "out", 0 0, L_0x5c7c3312bb10;  alias, 1 drivers
S_0x5c7c32d5bef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d5bcd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312bb10 .functor NAND 1, L_0x5c7c3312b250, L_0x5c7c3312b250, C4<1>, C4<1>;
v0x5c7c32d5c160_0 .net "in_a", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d5c220_0 .net "in_b", 0 0, L_0x5c7c3312b250;  alias, 1 drivers
v0x5c7c32d5c2e0_0 .net "out", 0 0, L_0x5c7c3312bb10;  alias, 1 drivers
S_0x5c7c32d5c5b0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d58810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d61ff0_0 .net "branch1_out", 0 0, L_0x5c7c3312be80;  1 drivers
v0x5c7c32d62120_0 .net "branch2_out", 0 0, L_0x5c7c3312c000;  1 drivers
v0x5c7c32d62270_0 .net "in_a", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
v0x5c7c32d62340_0 .net "in_b", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
v0x5c7c32d623e0_0 .net "out", 0 0, L_0x5c7c3312c180;  alias, 1 drivers
v0x5c7c32d62480_0 .net "temp1_out", 0 0, L_0x5c7c3312bdd0;  1 drivers
v0x5c7c32d62520_0 .net "temp2_out", 0 0, L_0x5c7c3312bf50;  1 drivers
v0x5c7c32d625c0_0 .net "temp3_out", 0 0, L_0x5c7c3312c0d0;  1 drivers
S_0x5c7c32d5c830 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d5c5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d5d830_0 .net "in_a", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
v0x5c7c32d5d8d0_0 .net "in_b", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
v0x5c7c32d5d990_0 .net "out", 0 0, L_0x5c7c3312bdd0;  alias, 1 drivers
v0x5c7c32d5dab0_0 .net "temp_out", 0 0, L_0x5c7c3312bd20;  1 drivers
S_0x5c7c32d5caa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d5c830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312bd20 .functor NAND 1, L_0x5c7c3312ba60, L_0x5c7c3312ba60, C4<1>, C4<1>;
v0x5c7c32d5cd10_0 .net "in_a", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
v0x5c7c32d5cdd0_0 .net "in_b", 0 0, L_0x5c7c3312ba60;  alias, 1 drivers
v0x5c7c32d5ce90_0 .net "out", 0 0, L_0x5c7c3312bd20;  alias, 1 drivers
S_0x5c7c32d5cf90 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d5c830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d5d680_0 .net "in_a", 0 0, L_0x5c7c3312bd20;  alias, 1 drivers
v0x5c7c32d5d720_0 .net "out", 0 0, L_0x5c7c3312bdd0;  alias, 1 drivers
S_0x5c7c32d5d160 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d5cf90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312bdd0 .functor NAND 1, L_0x5c7c3312bd20, L_0x5c7c3312bd20, C4<1>, C4<1>;
v0x5c7c32d5d3d0_0 .net "in_a", 0 0, L_0x5c7c3312bd20;  alias, 1 drivers
v0x5c7c32d5d490_0 .net "in_b", 0 0, L_0x5c7c3312bd20;  alias, 1 drivers
v0x5c7c32d5d580_0 .net "out", 0 0, L_0x5c7c3312bdd0;  alias, 1 drivers
S_0x5c7c32d5dc20 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d5c5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d5ec50_0 .net "in_a", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
v0x5c7c32d5ecf0_0 .net "in_b", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
v0x5c7c32d5edb0_0 .net "out", 0 0, L_0x5c7c3312bf50;  alias, 1 drivers
v0x5c7c32d5eed0_0 .net "temp_out", 0 0, L_0x5c7c32d60a70;  1 drivers
S_0x5c7c32d5de00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d5dc20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d60a70 .functor NAND 1, L_0x5c7c3312bc70, L_0x5c7c3312bc70, C4<1>, C4<1>;
v0x5c7c32d5e070_0 .net "in_a", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
v0x5c7c32d5e130_0 .net "in_b", 0 0, L_0x5c7c3312bc70;  alias, 1 drivers
v0x5c7c32d5e280_0 .net "out", 0 0, L_0x5c7c32d60a70;  alias, 1 drivers
S_0x5c7c32d5e380 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d5dc20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d5eaa0_0 .net "in_a", 0 0, L_0x5c7c32d60a70;  alias, 1 drivers
v0x5c7c32d5eb40_0 .net "out", 0 0, L_0x5c7c3312bf50;  alias, 1 drivers
S_0x5c7c32d5e550 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d5e380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312bf50 .functor NAND 1, L_0x5c7c32d60a70, L_0x5c7c32d60a70, C4<1>, C4<1>;
v0x5c7c32d5e7c0_0 .net "in_a", 0 0, L_0x5c7c32d60a70;  alias, 1 drivers
v0x5c7c32d5e8b0_0 .net "in_b", 0 0, L_0x5c7c32d60a70;  alias, 1 drivers
v0x5c7c32d5e9a0_0 .net "out", 0 0, L_0x5c7c3312bf50;  alias, 1 drivers
S_0x5c7c32d5f040 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d5c5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d60080_0 .net "in_a", 0 0, L_0x5c7c3312be80;  alias, 1 drivers
v0x5c7c32d60150_0 .net "in_b", 0 0, L_0x5c7c3312c000;  alias, 1 drivers
v0x5c7c32d60220_0 .net "out", 0 0, L_0x5c7c3312c0d0;  alias, 1 drivers
v0x5c7c32d60340_0 .net "temp_out", 0 0, L_0x5c7c32d613e0;  1 drivers
S_0x5c7c32d5f220 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d5f040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d613e0 .functor NAND 1, L_0x5c7c3312be80, L_0x5c7c3312c000, C4<1>, C4<1>;
v0x5c7c32d5f470_0 .net "in_a", 0 0, L_0x5c7c3312be80;  alias, 1 drivers
v0x5c7c32d5f550_0 .net "in_b", 0 0, L_0x5c7c3312c000;  alias, 1 drivers
v0x5c7c32d5f610_0 .net "out", 0 0, L_0x5c7c32d613e0;  alias, 1 drivers
S_0x5c7c32d5f760 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d5f040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d5fed0_0 .net "in_a", 0 0, L_0x5c7c32d613e0;  alias, 1 drivers
v0x5c7c32d5ff70_0 .net "out", 0 0, L_0x5c7c3312c0d0;  alias, 1 drivers
S_0x5c7c32d5f980 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d5f760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c0d0 .functor NAND 1, L_0x5c7c32d613e0, L_0x5c7c32d613e0, C4<1>, C4<1>;
v0x5c7c32d5fbf0_0 .net "in_a", 0 0, L_0x5c7c32d613e0;  alias, 1 drivers
v0x5c7c32d5fce0_0 .net "in_b", 0 0, L_0x5c7c32d613e0;  alias, 1 drivers
v0x5c7c32d5fdd0_0 .net "out", 0 0, L_0x5c7c3312c0d0;  alias, 1 drivers
S_0x5c7c32d60490 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d5c5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d60bc0_0 .net "in_a", 0 0, L_0x5c7c3312bdd0;  alias, 1 drivers
v0x5c7c32d60c60_0 .net "out", 0 0, L_0x5c7c3312be80;  alias, 1 drivers
S_0x5c7c32d60660 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d60490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312be80 .functor NAND 1, L_0x5c7c3312bdd0, L_0x5c7c3312bdd0, C4<1>, C4<1>;
v0x5c7c32d608d0_0 .net "in_a", 0 0, L_0x5c7c3312bdd0;  alias, 1 drivers
v0x5c7c32d60990_0 .net "in_b", 0 0, L_0x5c7c3312bdd0;  alias, 1 drivers
v0x5c7c32d60ae0_0 .net "out", 0 0, L_0x5c7c3312be80;  alias, 1 drivers
S_0x5c7c32d60d60 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d5c5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d61530_0 .net "in_a", 0 0, L_0x5c7c3312bf50;  alias, 1 drivers
v0x5c7c32d615d0_0 .net "out", 0 0, L_0x5c7c3312c000;  alias, 1 drivers
S_0x5c7c32d60fd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d60d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c000 .functor NAND 1, L_0x5c7c3312bf50, L_0x5c7c3312bf50, C4<1>, C4<1>;
v0x5c7c32d61240_0 .net "in_a", 0 0, L_0x5c7c3312bf50;  alias, 1 drivers
v0x5c7c32d61300_0 .net "in_b", 0 0, L_0x5c7c3312bf50;  alias, 1 drivers
v0x5c7c32d61450_0 .net "out", 0 0, L_0x5c7c3312c000;  alias, 1 drivers
S_0x5c7c32d616d0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d5c5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d61e70_0 .net "in_a", 0 0, L_0x5c7c3312c0d0;  alias, 1 drivers
v0x5c7c32d61f10_0 .net "out", 0 0, L_0x5c7c3312c180;  alias, 1 drivers
S_0x5c7c32d618f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d616d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c180 .functor NAND 1, L_0x5c7c3312c0d0, L_0x5c7c3312c0d0, C4<1>, C4<1>;
v0x5c7c32d61b60_0 .net "in_a", 0 0, L_0x5c7c3312c0d0;  alias, 1 drivers
v0x5c7c32d61c20_0 .net "in_b", 0 0, L_0x5c7c3312c0d0;  alias, 1 drivers
v0x5c7c32d61d70_0 .net "out", 0 0, L_0x5c7c3312c180;  alias, 1 drivers
S_0x5c7c32d630f0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32d4b0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d68ae0_0 .net "branch1_out", 0 0, L_0x5c7c3312c410;  1 drivers
v0x5c7c32d68c10_0 .net "branch2_out", 0 0, L_0x5c7c3312c6a0;  1 drivers
v0x5c7c32d68d60_0 .net "in_a", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d68f40_0 .net "in_b", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d690f0_0 .net "out", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d69190_0 .net "temp1_out", 0 0, L_0x5c7c3312c360;  1 drivers
v0x5c7c32d69230_0 .net "temp2_out", 0 0, L_0x5c7c3312c5f0;  1 drivers
v0x5c7c32d692d0_0 .net "temp3_out", 0 0, L_0x5c7c3312c880;  1 drivers
S_0x5c7c32d63280 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d630f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d64320_0 .net "in_a", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d643c0_0 .net "in_b", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d64480_0 .net "out", 0 0, L_0x5c7c3312c360;  alias, 1 drivers
v0x5c7c32d645a0_0 .net "temp_out", 0 0, L_0x5c7c32d61d00;  1 drivers
S_0x5c7c32d634a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d63280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d61d00 .functor NAND 1, L_0x5c7c3312a700, L_0x5c7c3312a700, C4<1>, C4<1>;
v0x5c7c32d63710_0 .net "in_a", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d63860_0 .net "in_b", 0 0, L_0x5c7c3312a700;  alias, 1 drivers
v0x5c7c32d63920_0 .net "out", 0 0, L_0x5c7c32d61d00;  alias, 1 drivers
S_0x5c7c32d63a50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d63280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d64170_0 .net "in_a", 0 0, L_0x5c7c32d61d00;  alias, 1 drivers
v0x5c7c32d64210_0 .net "out", 0 0, L_0x5c7c3312c360;  alias, 1 drivers
S_0x5c7c32d63c20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d63a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c360 .functor NAND 1, L_0x5c7c32d61d00, L_0x5c7c32d61d00, C4<1>, C4<1>;
v0x5c7c32d63e90_0 .net "in_a", 0 0, L_0x5c7c32d61d00;  alias, 1 drivers
v0x5c7c32d63f80_0 .net "in_b", 0 0, L_0x5c7c32d61d00;  alias, 1 drivers
v0x5c7c32d64070_0 .net "out", 0 0, L_0x5c7c3312c360;  alias, 1 drivers
S_0x5c7c32d64710 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d630f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d65740_0 .net "in_a", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d657e0_0 .net "in_b", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d658a0_0 .net "out", 0 0, L_0x5c7c3312c5f0;  alias, 1 drivers
v0x5c7c32d659c0_0 .net "temp_out", 0 0, L_0x5c7c32d67560;  1 drivers
S_0x5c7c32d648f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d64710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d67560 .functor NAND 1, L_0x5c7c3312b850, L_0x5c7c3312b850, C4<1>, C4<1>;
v0x5c7c32d64b60_0 .net "in_a", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d64cb0_0 .net "in_b", 0 0, L_0x5c7c3312b850;  alias, 1 drivers
v0x5c7c32d64d70_0 .net "out", 0 0, L_0x5c7c32d67560;  alias, 1 drivers
S_0x5c7c32d64e70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d64710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d65590_0 .net "in_a", 0 0, L_0x5c7c32d67560;  alias, 1 drivers
v0x5c7c32d65630_0 .net "out", 0 0, L_0x5c7c3312c5f0;  alias, 1 drivers
S_0x5c7c32d65040 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d64e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c5f0 .functor NAND 1, L_0x5c7c32d67560, L_0x5c7c32d67560, C4<1>, C4<1>;
v0x5c7c32d652b0_0 .net "in_a", 0 0, L_0x5c7c32d67560;  alias, 1 drivers
v0x5c7c32d653a0_0 .net "in_b", 0 0, L_0x5c7c32d67560;  alias, 1 drivers
v0x5c7c32d65490_0 .net "out", 0 0, L_0x5c7c3312c5f0;  alias, 1 drivers
S_0x5c7c32d65b30 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d630f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d66b70_0 .net "in_a", 0 0, L_0x5c7c3312c410;  alias, 1 drivers
v0x5c7c32d66c40_0 .net "in_b", 0 0, L_0x5c7c3312c6a0;  alias, 1 drivers
v0x5c7c32d66d10_0 .net "out", 0 0, L_0x5c7c3312c880;  alias, 1 drivers
v0x5c7c32d66e30_0 .net "temp_out", 0 0, L_0x5c7c32d67ed0;  1 drivers
S_0x5c7c32d65d10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d65b30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d67ed0 .functor NAND 1, L_0x5c7c3312c410, L_0x5c7c3312c6a0, C4<1>, C4<1>;
v0x5c7c32d65f60_0 .net "in_a", 0 0, L_0x5c7c3312c410;  alias, 1 drivers
v0x5c7c32d66040_0 .net "in_b", 0 0, L_0x5c7c3312c6a0;  alias, 1 drivers
v0x5c7c32d66100_0 .net "out", 0 0, L_0x5c7c32d67ed0;  alias, 1 drivers
S_0x5c7c32d66250 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d65b30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d669c0_0 .net "in_a", 0 0, L_0x5c7c32d67ed0;  alias, 1 drivers
v0x5c7c32d66a60_0 .net "out", 0 0, L_0x5c7c3312c880;  alias, 1 drivers
S_0x5c7c32d66470 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d66250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c880 .functor NAND 1, L_0x5c7c32d67ed0, L_0x5c7c32d67ed0, C4<1>, C4<1>;
v0x5c7c32d666e0_0 .net "in_a", 0 0, L_0x5c7c32d67ed0;  alias, 1 drivers
v0x5c7c32d667d0_0 .net "in_b", 0 0, L_0x5c7c32d67ed0;  alias, 1 drivers
v0x5c7c32d668c0_0 .net "out", 0 0, L_0x5c7c3312c880;  alias, 1 drivers
S_0x5c7c32d66f80 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d630f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d676b0_0 .net "in_a", 0 0, L_0x5c7c3312c360;  alias, 1 drivers
v0x5c7c32d67750_0 .net "out", 0 0, L_0x5c7c3312c410;  alias, 1 drivers
S_0x5c7c32d67150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d66f80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c410 .functor NAND 1, L_0x5c7c3312c360, L_0x5c7c3312c360, C4<1>, C4<1>;
v0x5c7c32d673c0_0 .net "in_a", 0 0, L_0x5c7c3312c360;  alias, 1 drivers
v0x5c7c32d67480_0 .net "in_b", 0 0, L_0x5c7c3312c360;  alias, 1 drivers
v0x5c7c32d675d0_0 .net "out", 0 0, L_0x5c7c3312c410;  alias, 1 drivers
S_0x5c7c32d67850 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d630f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d68020_0 .net "in_a", 0 0, L_0x5c7c3312c5f0;  alias, 1 drivers
v0x5c7c32d680c0_0 .net "out", 0 0, L_0x5c7c3312c6a0;  alias, 1 drivers
S_0x5c7c32d67ac0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d67850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c6a0 .functor NAND 1, L_0x5c7c3312c5f0, L_0x5c7c3312c5f0, C4<1>, C4<1>;
v0x5c7c32d67d30_0 .net "in_a", 0 0, L_0x5c7c3312c5f0;  alias, 1 drivers
v0x5c7c32d67df0_0 .net "in_b", 0 0, L_0x5c7c3312c5f0;  alias, 1 drivers
v0x5c7c32d67f40_0 .net "out", 0 0, L_0x5c7c3312c6a0;  alias, 1 drivers
S_0x5c7c32d681c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d630f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d68960_0 .net "in_a", 0 0, L_0x5c7c3312c880;  alias, 1 drivers
v0x5c7c32d68a00_0 .net "out", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
S_0x5c7c32d683e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d681c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312c930 .functor NAND 1, L_0x5c7c3312c880, L_0x5c7c3312c880, C4<1>, C4<1>;
v0x5c7c32d68650_0 .net "in_a", 0 0, L_0x5c7c3312c880;  alias, 1 drivers
v0x5c7c32d68710_0 .net "in_b", 0 0, L_0x5c7c3312c880;  alias, 1 drivers
v0x5c7c32d68860_0 .net "out", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
S_0x5c7c32d69930 .scope module, "fa_gate13" "FullAdder" 2 18, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32d87c00_0 .net "a", 0 0, L_0x5c7c3312f0f0;  1 drivers
v0x5c7c32d87ca0_0 .net "b", 0 0, L_0x5c7c3312f190;  1 drivers
v0x5c7c32d87d60_0 .net "c", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d87e00_0 .net "carry", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d87ea0_0 .net "sum", 0 0, L_0x5c7c3312e7a0;  1 drivers
v0x5c7c32d87f40_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c3312cd20;  1 drivers
v0x5c7c32d87fe0_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c3312de70;  1 drivers
v0x5c7c32d88080_0 .net "tmp_sum_out", 0 0, L_0x5c7c3312d870;  1 drivers
S_0x5c7c32d69b10 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32d69930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d75620_0 .net "a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d757d0_0 .net "b", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d759a0_0 .net "carry", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d75a40_0 .net "sum", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
S_0x5c7c32d69d10 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d69b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d6ae00_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6aed0_0 .net "in_b", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6afa0_0 .net "out", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d6b0c0_0 .net "temp_out", 0 0, L_0x5c7c32d687f0;  1 drivers
S_0x5c7c32d69f80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d69d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d687f0 .functor NAND 1, L_0x5c7c3312f0f0, L_0x5c7c3312f190, C4<1>, C4<1>;
v0x5c7c32d6a1f0_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6a2d0_0 .net "in_b", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6a390_0 .net "out", 0 0, L_0x5c7c32d687f0;  alias, 1 drivers
S_0x5c7c32d6a4e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d69d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d6ac50_0 .net "in_a", 0 0, L_0x5c7c32d687f0;  alias, 1 drivers
v0x5c7c32d6acf0_0 .net "out", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
S_0x5c7c32d6a700 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d6a4e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312cd20 .functor NAND 1, L_0x5c7c32d687f0, L_0x5c7c32d687f0, C4<1>, C4<1>;
v0x5c7c32d6a970_0 .net "in_a", 0 0, L_0x5c7c32d687f0;  alias, 1 drivers
v0x5c7c32d6aa60_0 .net "in_b", 0 0, L_0x5c7c32d687f0;  alias, 1 drivers
v0x5c7c32d6ab50_0 .net "out", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
S_0x5c7c32d6b180 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d69b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d74f40_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d74fe0_0 .net "in_b", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d750a0_0 .net "out", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d75140_0 .net "temp_a_and_out", 0 0, L_0x5c7c3312cf30;  1 drivers
v0x5c7c32d752f0_0 .net "temp_a_out", 0 0, L_0x5c7c3312cdd0;  1 drivers
v0x5c7c32d75390_0 .net "temp_b_and_out", 0 0, L_0x5c7c3312d140;  1 drivers
v0x5c7c32d75540_0 .net "temp_b_out", 0 0, L_0x5c7c3312cfe0;  1 drivers
S_0x5c7c32d6b360 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d6b180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d6c420_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6c4c0_0 .net "in_b", 0 0, L_0x5c7c3312cdd0;  alias, 1 drivers
v0x5c7c32d6c5b0_0 .net "out", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
v0x5c7c32d6c6d0_0 .net "temp_out", 0 0, L_0x5c7c3312ce80;  1 drivers
S_0x5c7c32d6b5d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d6b360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ce80 .functor NAND 1, L_0x5c7c3312f0f0, L_0x5c7c3312cdd0, C4<1>, C4<1>;
v0x5c7c32d6b840_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6b950_0 .net "in_b", 0 0, L_0x5c7c3312cdd0;  alias, 1 drivers
v0x5c7c32d6ba10_0 .net "out", 0 0, L_0x5c7c3312ce80;  alias, 1 drivers
S_0x5c7c32d6bb30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d6b360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d6c270_0 .net "in_a", 0 0, L_0x5c7c3312ce80;  alias, 1 drivers
v0x5c7c32d6c310_0 .net "out", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
S_0x5c7c32d6bd50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d6bb30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312cf30 .functor NAND 1, L_0x5c7c3312ce80, L_0x5c7c3312ce80, C4<1>, C4<1>;
v0x5c7c32d6bfc0_0 .net "in_a", 0 0, L_0x5c7c3312ce80;  alias, 1 drivers
v0x5c7c32d6c080_0 .net "in_b", 0 0, L_0x5c7c3312ce80;  alias, 1 drivers
v0x5c7c32d6c170_0 .net "out", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
S_0x5c7c32d6c790 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d6b180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d6d7c0_0 .net "in_a", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6d860_0 .net "in_b", 0 0, L_0x5c7c3312cfe0;  alias, 1 drivers
v0x5c7c32d6d950_0 .net "out", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
v0x5c7c32d6da70_0 .net "temp_out", 0 0, L_0x5c7c3312d090;  1 drivers
S_0x5c7c32d6c970 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d6c790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d090 .functor NAND 1, L_0x5c7c3312f190, L_0x5c7c3312cfe0, C4<1>, C4<1>;
v0x5c7c32d6cbe0_0 .net "in_a", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6ccf0_0 .net "in_b", 0 0, L_0x5c7c3312cfe0;  alias, 1 drivers
v0x5c7c32d6cdb0_0 .net "out", 0 0, L_0x5c7c3312d090;  alias, 1 drivers
S_0x5c7c32d6ced0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d6c790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d6d610_0 .net "in_a", 0 0, L_0x5c7c3312d090;  alias, 1 drivers
v0x5c7c32d6d6b0_0 .net "out", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
S_0x5c7c32d6d0f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d6ced0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d140 .functor NAND 1, L_0x5c7c3312d090, L_0x5c7c3312d090, C4<1>, C4<1>;
v0x5c7c32d6d360_0 .net "in_a", 0 0, L_0x5c7c3312d090;  alias, 1 drivers
v0x5c7c32d6d420_0 .net "in_b", 0 0, L_0x5c7c3312d090;  alias, 1 drivers
v0x5c7c32d6d510_0 .net "out", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
S_0x5c7c32d6dbc0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d6b180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d6e300_0 .net "in_a", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6e3a0_0 .net "out", 0 0, L_0x5c7c3312cdd0;  alias, 1 drivers
S_0x5c7c32d6dd90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d6dbc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312cdd0 .functor NAND 1, L_0x5c7c3312f190, L_0x5c7c3312f190, C4<1>, C4<1>;
v0x5c7c32d6dfe0_0 .net "in_a", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6e130_0 .net "in_b", 0 0, L_0x5c7c3312f190;  alias, 1 drivers
v0x5c7c32d6e1f0_0 .net "out", 0 0, L_0x5c7c3312cdd0;  alias, 1 drivers
S_0x5c7c32d6e4a0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d6b180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d6ec20_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6ecc0_0 .net "out", 0 0, L_0x5c7c3312cfe0;  alias, 1 drivers
S_0x5c7c32d6e6c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d6e4a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312cfe0 .functor NAND 1, L_0x5c7c3312f0f0, L_0x5c7c3312f0f0, C4<1>, C4<1>;
v0x5c7c32d6e930_0 .net "in_a", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6ea80_0 .net "in_b", 0 0, L_0x5c7c3312f0f0;  alias, 1 drivers
v0x5c7c32d6eb40_0 .net "out", 0 0, L_0x5c7c3312cfe0;  alias, 1 drivers
S_0x5c7c32d6edc0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d6b180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d74890_0 .net "branch1_out", 0 0, L_0x5c7c3312d350;  1 drivers
v0x5c7c32d749c0_0 .net "branch2_out", 0 0, L_0x5c7c3312d5e0;  1 drivers
v0x5c7c32d74b10_0 .net "in_a", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
v0x5c7c32d74be0_0 .net "in_b", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
v0x5c7c32d74c80_0 .net "out", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d74d20_0 .net "temp1_out", 0 0, L_0x5c7c3312d2a0;  1 drivers
v0x5c7c32d74dc0_0 .net "temp2_out", 0 0, L_0x5c7c3312d530;  1 drivers
v0x5c7c32d74e60_0 .net "temp3_out", 0 0, L_0x5c7c3312d7c0;  1 drivers
S_0x5c7c32d6f040 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d6edc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d700d0_0 .net "in_a", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
v0x5c7c32d70170_0 .net "in_b", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
v0x5c7c32d70230_0 .net "out", 0 0, L_0x5c7c3312d2a0;  alias, 1 drivers
v0x5c7c32d70350_0 .net "temp_out", 0 0, L_0x5c7c3312d1f0;  1 drivers
S_0x5c7c32d6f2b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d6f040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d1f0 .functor NAND 1, L_0x5c7c3312cf30, L_0x5c7c3312cf30, C4<1>, C4<1>;
v0x5c7c32d6f520_0 .net "in_a", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
v0x5c7c32d6f5e0_0 .net "in_b", 0 0, L_0x5c7c3312cf30;  alias, 1 drivers
v0x5c7c32d6f730_0 .net "out", 0 0, L_0x5c7c3312d1f0;  alias, 1 drivers
S_0x5c7c32d6f830 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d6f040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d6ff20_0 .net "in_a", 0 0, L_0x5c7c3312d1f0;  alias, 1 drivers
v0x5c7c32d6ffc0_0 .net "out", 0 0, L_0x5c7c3312d2a0;  alias, 1 drivers
S_0x5c7c32d6fa00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d6f830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d2a0 .functor NAND 1, L_0x5c7c3312d1f0, L_0x5c7c3312d1f0, C4<1>, C4<1>;
v0x5c7c32d6fc70_0 .net "in_a", 0 0, L_0x5c7c3312d1f0;  alias, 1 drivers
v0x5c7c32d6fd30_0 .net "in_b", 0 0, L_0x5c7c3312d1f0;  alias, 1 drivers
v0x5c7c32d6fe20_0 .net "out", 0 0, L_0x5c7c3312d2a0;  alias, 1 drivers
S_0x5c7c32d704c0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d6edc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d714f0_0 .net "in_a", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
v0x5c7c32d71590_0 .net "in_b", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
v0x5c7c32d71650_0 .net "out", 0 0, L_0x5c7c3312d530;  alias, 1 drivers
v0x5c7c32d71770_0 .net "temp_out", 0 0, L_0x5c7c32d73310;  1 drivers
S_0x5c7c32d706a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d704c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d73310 .functor NAND 1, L_0x5c7c3312d140, L_0x5c7c3312d140, C4<1>, C4<1>;
v0x5c7c32d70910_0 .net "in_a", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
v0x5c7c32d709d0_0 .net "in_b", 0 0, L_0x5c7c3312d140;  alias, 1 drivers
v0x5c7c32d70b20_0 .net "out", 0 0, L_0x5c7c32d73310;  alias, 1 drivers
S_0x5c7c32d70c20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d704c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d71340_0 .net "in_a", 0 0, L_0x5c7c32d73310;  alias, 1 drivers
v0x5c7c32d713e0_0 .net "out", 0 0, L_0x5c7c3312d530;  alias, 1 drivers
S_0x5c7c32d70df0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d70c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d530 .functor NAND 1, L_0x5c7c32d73310, L_0x5c7c32d73310, C4<1>, C4<1>;
v0x5c7c32d71060_0 .net "in_a", 0 0, L_0x5c7c32d73310;  alias, 1 drivers
v0x5c7c32d71150_0 .net "in_b", 0 0, L_0x5c7c32d73310;  alias, 1 drivers
v0x5c7c32d71240_0 .net "out", 0 0, L_0x5c7c3312d530;  alias, 1 drivers
S_0x5c7c32d718e0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d6edc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d72920_0 .net "in_a", 0 0, L_0x5c7c3312d350;  alias, 1 drivers
v0x5c7c32d729f0_0 .net "in_b", 0 0, L_0x5c7c3312d5e0;  alias, 1 drivers
v0x5c7c32d72ac0_0 .net "out", 0 0, L_0x5c7c3312d7c0;  alias, 1 drivers
v0x5c7c32d72be0_0 .net "temp_out", 0 0, L_0x5c7c32d73c80;  1 drivers
S_0x5c7c32d71ac0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d718e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d73c80 .functor NAND 1, L_0x5c7c3312d350, L_0x5c7c3312d5e0, C4<1>, C4<1>;
v0x5c7c32d71d10_0 .net "in_a", 0 0, L_0x5c7c3312d350;  alias, 1 drivers
v0x5c7c32d71df0_0 .net "in_b", 0 0, L_0x5c7c3312d5e0;  alias, 1 drivers
v0x5c7c32d71eb0_0 .net "out", 0 0, L_0x5c7c32d73c80;  alias, 1 drivers
S_0x5c7c32d72000 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d718e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d72770_0 .net "in_a", 0 0, L_0x5c7c32d73c80;  alias, 1 drivers
v0x5c7c32d72810_0 .net "out", 0 0, L_0x5c7c3312d7c0;  alias, 1 drivers
S_0x5c7c32d72220 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d72000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d7c0 .functor NAND 1, L_0x5c7c32d73c80, L_0x5c7c32d73c80, C4<1>, C4<1>;
v0x5c7c32d72490_0 .net "in_a", 0 0, L_0x5c7c32d73c80;  alias, 1 drivers
v0x5c7c32d72580_0 .net "in_b", 0 0, L_0x5c7c32d73c80;  alias, 1 drivers
v0x5c7c32d72670_0 .net "out", 0 0, L_0x5c7c3312d7c0;  alias, 1 drivers
S_0x5c7c32d72d30 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d6edc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d73460_0 .net "in_a", 0 0, L_0x5c7c3312d2a0;  alias, 1 drivers
v0x5c7c32d73500_0 .net "out", 0 0, L_0x5c7c3312d350;  alias, 1 drivers
S_0x5c7c32d72f00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d72d30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d350 .functor NAND 1, L_0x5c7c3312d2a0, L_0x5c7c3312d2a0, C4<1>, C4<1>;
v0x5c7c32d73170_0 .net "in_a", 0 0, L_0x5c7c3312d2a0;  alias, 1 drivers
v0x5c7c32d73230_0 .net "in_b", 0 0, L_0x5c7c3312d2a0;  alias, 1 drivers
v0x5c7c32d73380_0 .net "out", 0 0, L_0x5c7c3312d350;  alias, 1 drivers
S_0x5c7c32d73600 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d6edc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d73dd0_0 .net "in_a", 0 0, L_0x5c7c3312d530;  alias, 1 drivers
v0x5c7c32d73e70_0 .net "out", 0 0, L_0x5c7c3312d5e0;  alias, 1 drivers
S_0x5c7c32d73870 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d73600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d5e0 .functor NAND 1, L_0x5c7c3312d530, L_0x5c7c3312d530, C4<1>, C4<1>;
v0x5c7c32d73ae0_0 .net "in_a", 0 0, L_0x5c7c3312d530;  alias, 1 drivers
v0x5c7c32d73ba0_0 .net "in_b", 0 0, L_0x5c7c3312d530;  alias, 1 drivers
v0x5c7c32d73cf0_0 .net "out", 0 0, L_0x5c7c3312d5e0;  alias, 1 drivers
S_0x5c7c32d73f70 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d6edc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d74710_0 .net "in_a", 0 0, L_0x5c7c3312d7c0;  alias, 1 drivers
v0x5c7c32d747b0_0 .net "out", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
S_0x5c7c32d74190 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d73f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312d870 .functor NAND 1, L_0x5c7c3312d7c0, L_0x5c7c3312d7c0, C4<1>, C4<1>;
v0x5c7c32d74400_0 .net "in_a", 0 0, L_0x5c7c3312d7c0;  alias, 1 drivers
v0x5c7c32d744c0_0 .net "in_b", 0 0, L_0x5c7c3312d7c0;  alias, 1 drivers
v0x5c7c32d74610_0 .net "out", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
S_0x5c7c32d75b20 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32d69930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d815d0_0 .net "a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d81670_0 .net "b", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d81730_0 .net "carry", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d817d0_0 .net "sum", 0 0, L_0x5c7c3312e7a0;  alias, 1 drivers
S_0x5c7c32d75cd0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d75b20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d76c70_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d76d10_0 .net "in_b", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d76dd0_0 .net "out", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d76ef0_0 .net "temp_out", 0 0, L_0x5c7c32d745a0;  1 drivers
S_0x5c7c32d75e80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d75cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d745a0 .functor NAND 1, L_0x5c7c3312d870, L_0x5c7c3312c930, C4<1>, C4<1>;
v0x5c7c32d760f0_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d761b0_0 .net "in_b", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d76270_0 .net "out", 0 0, L_0x5c7c32d745a0;  alias, 1 drivers
S_0x5c7c32d763a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d75cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d76ac0_0 .net "in_a", 0 0, L_0x5c7c32d745a0;  alias, 1 drivers
v0x5c7c32d76b60_0 .net "out", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
S_0x5c7c32d76570 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d763a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312de70 .functor NAND 1, L_0x5c7c32d745a0, L_0x5c7c32d745a0, C4<1>, C4<1>;
v0x5c7c32d767e0_0 .net "in_a", 0 0, L_0x5c7c32d745a0;  alias, 1 drivers
v0x5c7c32d768d0_0 .net "in_b", 0 0, L_0x5c7c32d745a0;  alias, 1 drivers
v0x5c7c32d769c0_0 .net "out", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
S_0x5c7c32d77060 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d75b20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d80ef0_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d80f90_0 .net "in_b", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d81050_0 .net "out", 0 0, L_0x5c7c3312e7a0;  alias, 1 drivers
v0x5c7c32d810f0_0 .net "temp_a_and_out", 0 0, L_0x5c7c3312e080;  1 drivers
v0x5c7c32d812a0_0 .net "temp_a_out", 0 0, L_0x5c7c3312df20;  1 drivers
v0x5c7c32d81340_0 .net "temp_b_and_out", 0 0, L_0x5c7c3312e290;  1 drivers
v0x5c7c32d814f0_0 .net "temp_b_out", 0 0, L_0x5c7c3312e130;  1 drivers
S_0x5c7c32d77240 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d77060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d782e0_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d78490_0 .net "in_b", 0 0, L_0x5c7c3312df20;  alias, 1 drivers
v0x5c7c32d78580_0 .net "out", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
v0x5c7c32d786a0_0 .net "temp_out", 0 0, L_0x5c7c3312dfd0;  1 drivers
S_0x5c7c32d774b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d77240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312dfd0 .functor NAND 1, L_0x5c7c3312d870, L_0x5c7c3312df20, C4<1>, C4<1>;
v0x5c7c32d77720_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d777e0_0 .net "in_b", 0 0, L_0x5c7c3312df20;  alias, 1 drivers
v0x5c7c32d778a0_0 .net "out", 0 0, L_0x5c7c3312dfd0;  alias, 1 drivers
S_0x5c7c32d779c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d77240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d78130_0 .net "in_a", 0 0, L_0x5c7c3312dfd0;  alias, 1 drivers
v0x5c7c32d781d0_0 .net "out", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
S_0x5c7c32d77be0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d779c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e080 .functor NAND 1, L_0x5c7c3312dfd0, L_0x5c7c3312dfd0, C4<1>, C4<1>;
v0x5c7c32d77e50_0 .net "in_a", 0 0, L_0x5c7c3312dfd0;  alias, 1 drivers
v0x5c7c32d77f40_0 .net "in_b", 0 0, L_0x5c7c3312dfd0;  alias, 1 drivers
v0x5c7c32d78030_0 .net "out", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
S_0x5c7c32d78760 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d77060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d79770_0 .net "in_a", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d79810_0 .net "in_b", 0 0, L_0x5c7c3312e130;  alias, 1 drivers
v0x5c7c32d79900_0 .net "out", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
v0x5c7c32d79a20_0 .net "temp_out", 0 0, L_0x5c7c3312e1e0;  1 drivers
S_0x5c7c32d78940 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d78760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e1e0 .functor NAND 1, L_0x5c7c3312c930, L_0x5c7c3312e130, C4<1>, C4<1>;
v0x5c7c32d78bb0_0 .net "in_a", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d78c70_0 .net "in_b", 0 0, L_0x5c7c3312e130;  alias, 1 drivers
v0x5c7c32d78d30_0 .net "out", 0 0, L_0x5c7c3312e1e0;  alias, 1 drivers
S_0x5c7c32d78e50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d78760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d795c0_0 .net "in_a", 0 0, L_0x5c7c3312e1e0;  alias, 1 drivers
v0x5c7c32d79660_0 .net "out", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
S_0x5c7c32d79070 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d78e50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e290 .functor NAND 1, L_0x5c7c3312e1e0, L_0x5c7c3312e1e0, C4<1>, C4<1>;
v0x5c7c32d792e0_0 .net "in_a", 0 0, L_0x5c7c3312e1e0;  alias, 1 drivers
v0x5c7c32d793d0_0 .net "in_b", 0 0, L_0x5c7c3312e1e0;  alias, 1 drivers
v0x5c7c32d794c0_0 .net "out", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
S_0x5c7c32d79b70 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d77060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7a380_0 .net "in_a", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d7a420_0 .net "out", 0 0, L_0x5c7c3312df20;  alias, 1 drivers
S_0x5c7c32d79d40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d79b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312df20 .functor NAND 1, L_0x5c7c3312c930, L_0x5c7c3312c930, C4<1>, C4<1>;
v0x5c7c32d79f90_0 .net "in_a", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d7a160_0 .net "in_b", 0 0, L_0x5c7c3312c930;  alias, 1 drivers
v0x5c7c32d7a220_0 .net "out", 0 0, L_0x5c7c3312df20;  alias, 1 drivers
S_0x5c7c32d7a520 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d77060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7ac60_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d7ad00_0 .net "out", 0 0, L_0x5c7c3312e130;  alias, 1 drivers
S_0x5c7c32d7a740 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7a520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e130 .functor NAND 1, L_0x5c7c3312d870, L_0x5c7c3312d870, C4<1>, C4<1>;
v0x5c7c32d7a9b0_0 .net "in_a", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d7aa70_0 .net "in_b", 0 0, L_0x5c7c3312d870;  alias, 1 drivers
v0x5c7c32d7ab30_0 .net "out", 0 0, L_0x5c7c3312e130;  alias, 1 drivers
S_0x5c7c32d7ae00 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d77060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d80840_0 .net "branch1_out", 0 0, L_0x5c7c3312e4a0;  1 drivers
v0x5c7c32d80970_0 .net "branch2_out", 0 0, L_0x5c7c3312e620;  1 drivers
v0x5c7c32d80ac0_0 .net "in_a", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
v0x5c7c32d80b90_0 .net "in_b", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
v0x5c7c32d80c30_0 .net "out", 0 0, L_0x5c7c3312e7a0;  alias, 1 drivers
v0x5c7c32d80cd0_0 .net "temp1_out", 0 0, L_0x5c7c3312e3f0;  1 drivers
v0x5c7c32d80d70_0 .net "temp2_out", 0 0, L_0x5c7c3312e570;  1 drivers
v0x5c7c32d80e10_0 .net "temp3_out", 0 0, L_0x5c7c3312e6f0;  1 drivers
S_0x5c7c32d7b080 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d7ae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d7c080_0 .net "in_a", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
v0x5c7c32d7c120_0 .net "in_b", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
v0x5c7c32d7c1e0_0 .net "out", 0 0, L_0x5c7c3312e3f0;  alias, 1 drivers
v0x5c7c32d7c300_0 .net "temp_out", 0 0, L_0x5c7c3312e340;  1 drivers
S_0x5c7c32d7b2f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d7b080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e340 .functor NAND 1, L_0x5c7c3312e080, L_0x5c7c3312e080, C4<1>, C4<1>;
v0x5c7c32d7b560_0 .net "in_a", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
v0x5c7c32d7b620_0 .net "in_b", 0 0, L_0x5c7c3312e080;  alias, 1 drivers
v0x5c7c32d7b6e0_0 .net "out", 0 0, L_0x5c7c3312e340;  alias, 1 drivers
S_0x5c7c32d7b7e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d7b080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7bed0_0 .net "in_a", 0 0, L_0x5c7c3312e340;  alias, 1 drivers
v0x5c7c32d7bf70_0 .net "out", 0 0, L_0x5c7c3312e3f0;  alias, 1 drivers
S_0x5c7c32d7b9b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7b7e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e3f0 .functor NAND 1, L_0x5c7c3312e340, L_0x5c7c3312e340, C4<1>, C4<1>;
v0x5c7c32d7bc20_0 .net "in_a", 0 0, L_0x5c7c3312e340;  alias, 1 drivers
v0x5c7c32d7bce0_0 .net "in_b", 0 0, L_0x5c7c3312e340;  alias, 1 drivers
v0x5c7c32d7bdd0_0 .net "out", 0 0, L_0x5c7c3312e3f0;  alias, 1 drivers
S_0x5c7c32d7c470 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d7ae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d7d4a0_0 .net "in_a", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
v0x5c7c32d7d540_0 .net "in_b", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
v0x5c7c32d7d600_0 .net "out", 0 0, L_0x5c7c3312e570;  alias, 1 drivers
v0x5c7c32d7d720_0 .net "temp_out", 0 0, L_0x5c7c32d7f2c0;  1 drivers
S_0x5c7c32d7c650 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d7c470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d7f2c0 .functor NAND 1, L_0x5c7c3312e290, L_0x5c7c3312e290, C4<1>, C4<1>;
v0x5c7c32d7c8c0_0 .net "in_a", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
v0x5c7c32d7c980_0 .net "in_b", 0 0, L_0x5c7c3312e290;  alias, 1 drivers
v0x5c7c32d7cad0_0 .net "out", 0 0, L_0x5c7c32d7f2c0;  alias, 1 drivers
S_0x5c7c32d7cbd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d7c470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7d2f0_0 .net "in_a", 0 0, L_0x5c7c32d7f2c0;  alias, 1 drivers
v0x5c7c32d7d390_0 .net "out", 0 0, L_0x5c7c3312e570;  alias, 1 drivers
S_0x5c7c32d7cda0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7cbd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e570 .functor NAND 1, L_0x5c7c32d7f2c0, L_0x5c7c32d7f2c0, C4<1>, C4<1>;
v0x5c7c32d7d010_0 .net "in_a", 0 0, L_0x5c7c32d7f2c0;  alias, 1 drivers
v0x5c7c32d7d100_0 .net "in_b", 0 0, L_0x5c7c32d7f2c0;  alias, 1 drivers
v0x5c7c32d7d1f0_0 .net "out", 0 0, L_0x5c7c3312e570;  alias, 1 drivers
S_0x5c7c32d7d890 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d7ae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d7e8d0_0 .net "in_a", 0 0, L_0x5c7c3312e4a0;  alias, 1 drivers
v0x5c7c32d7e9a0_0 .net "in_b", 0 0, L_0x5c7c3312e620;  alias, 1 drivers
v0x5c7c32d7ea70_0 .net "out", 0 0, L_0x5c7c3312e6f0;  alias, 1 drivers
v0x5c7c32d7eb90_0 .net "temp_out", 0 0, L_0x5c7c32d7fc30;  1 drivers
S_0x5c7c32d7da70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d7d890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d7fc30 .functor NAND 1, L_0x5c7c3312e4a0, L_0x5c7c3312e620, C4<1>, C4<1>;
v0x5c7c32d7dcc0_0 .net "in_a", 0 0, L_0x5c7c3312e4a0;  alias, 1 drivers
v0x5c7c32d7dda0_0 .net "in_b", 0 0, L_0x5c7c3312e620;  alias, 1 drivers
v0x5c7c32d7de60_0 .net "out", 0 0, L_0x5c7c32d7fc30;  alias, 1 drivers
S_0x5c7c32d7dfb0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d7d890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7e720_0 .net "in_a", 0 0, L_0x5c7c32d7fc30;  alias, 1 drivers
v0x5c7c32d7e7c0_0 .net "out", 0 0, L_0x5c7c3312e6f0;  alias, 1 drivers
S_0x5c7c32d7e1d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7dfb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e6f0 .functor NAND 1, L_0x5c7c32d7fc30, L_0x5c7c32d7fc30, C4<1>, C4<1>;
v0x5c7c32d7e440_0 .net "in_a", 0 0, L_0x5c7c32d7fc30;  alias, 1 drivers
v0x5c7c32d7e530_0 .net "in_b", 0 0, L_0x5c7c32d7fc30;  alias, 1 drivers
v0x5c7c32d7e620_0 .net "out", 0 0, L_0x5c7c3312e6f0;  alias, 1 drivers
S_0x5c7c32d7ece0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d7ae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7f410_0 .net "in_a", 0 0, L_0x5c7c3312e3f0;  alias, 1 drivers
v0x5c7c32d7f4b0_0 .net "out", 0 0, L_0x5c7c3312e4a0;  alias, 1 drivers
S_0x5c7c32d7eeb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7ece0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e4a0 .functor NAND 1, L_0x5c7c3312e3f0, L_0x5c7c3312e3f0, C4<1>, C4<1>;
v0x5c7c32d7f120_0 .net "in_a", 0 0, L_0x5c7c3312e3f0;  alias, 1 drivers
v0x5c7c32d7f1e0_0 .net "in_b", 0 0, L_0x5c7c3312e3f0;  alias, 1 drivers
v0x5c7c32d7f330_0 .net "out", 0 0, L_0x5c7c3312e4a0;  alias, 1 drivers
S_0x5c7c32d7f5b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d7ae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d7fd80_0 .net "in_a", 0 0, L_0x5c7c3312e570;  alias, 1 drivers
v0x5c7c32d7fe20_0 .net "out", 0 0, L_0x5c7c3312e620;  alias, 1 drivers
S_0x5c7c32d7f820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7f5b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e620 .functor NAND 1, L_0x5c7c3312e570, L_0x5c7c3312e570, C4<1>, C4<1>;
v0x5c7c32d7fa90_0 .net "in_a", 0 0, L_0x5c7c3312e570;  alias, 1 drivers
v0x5c7c32d7fb50_0 .net "in_b", 0 0, L_0x5c7c3312e570;  alias, 1 drivers
v0x5c7c32d7fca0_0 .net "out", 0 0, L_0x5c7c3312e620;  alias, 1 drivers
S_0x5c7c32d7ff20 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d7ae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d806c0_0 .net "in_a", 0 0, L_0x5c7c3312e6f0;  alias, 1 drivers
v0x5c7c32d80760_0 .net "out", 0 0, L_0x5c7c3312e7a0;  alias, 1 drivers
S_0x5c7c32d80140 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d7ff20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e7a0 .functor NAND 1, L_0x5c7c3312e6f0, L_0x5c7c3312e6f0, C4<1>, C4<1>;
v0x5c7c32d803b0_0 .net "in_a", 0 0, L_0x5c7c3312e6f0;  alias, 1 drivers
v0x5c7c32d80470_0 .net "in_b", 0 0, L_0x5c7c3312e6f0;  alias, 1 drivers
v0x5c7c32d805c0_0 .net "out", 0 0, L_0x5c7c3312e7a0;  alias, 1 drivers
S_0x5c7c32d81940 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32d69930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d87330_0 .net "branch1_out", 0 0, L_0x5c7c3312ea30;  1 drivers
v0x5c7c32d87460_0 .net "branch2_out", 0 0, L_0x5c7c3312ecc0;  1 drivers
v0x5c7c32d875b0_0 .net "in_a", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d87790_0 .net "in_b", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d87940_0 .net "out", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d879e0_0 .net "temp1_out", 0 0, L_0x5c7c3312e980;  1 drivers
v0x5c7c32d87a80_0 .net "temp2_out", 0 0, L_0x5c7c3312ec10;  1 drivers
v0x5c7c32d87b20_0 .net "temp3_out", 0 0, L_0x5c7c3312eea0;  1 drivers
S_0x5c7c32d81ad0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d81940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d82b70_0 .net "in_a", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d82c10_0 .net "in_b", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d82cd0_0 .net "out", 0 0, L_0x5c7c3312e980;  alias, 1 drivers
v0x5c7c32d82df0_0 .net "temp_out", 0 0, L_0x5c7c32d80550;  1 drivers
S_0x5c7c32d81cf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d81ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d80550 .functor NAND 1, L_0x5c7c3312cd20, L_0x5c7c3312cd20, C4<1>, C4<1>;
v0x5c7c32d81f60_0 .net "in_a", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d820b0_0 .net "in_b", 0 0, L_0x5c7c3312cd20;  alias, 1 drivers
v0x5c7c32d82170_0 .net "out", 0 0, L_0x5c7c32d80550;  alias, 1 drivers
S_0x5c7c32d822a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d81ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d829c0_0 .net "in_a", 0 0, L_0x5c7c32d80550;  alias, 1 drivers
v0x5c7c32d82a60_0 .net "out", 0 0, L_0x5c7c3312e980;  alias, 1 drivers
S_0x5c7c32d82470 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d822a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312e980 .functor NAND 1, L_0x5c7c32d80550, L_0x5c7c32d80550, C4<1>, C4<1>;
v0x5c7c32d826e0_0 .net "in_a", 0 0, L_0x5c7c32d80550;  alias, 1 drivers
v0x5c7c32d827d0_0 .net "in_b", 0 0, L_0x5c7c32d80550;  alias, 1 drivers
v0x5c7c32d828c0_0 .net "out", 0 0, L_0x5c7c3312e980;  alias, 1 drivers
S_0x5c7c32d82f60 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d81940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d83f90_0 .net "in_a", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d84030_0 .net "in_b", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d840f0_0 .net "out", 0 0, L_0x5c7c3312ec10;  alias, 1 drivers
v0x5c7c32d84210_0 .net "temp_out", 0 0, L_0x5c7c32d85db0;  1 drivers
S_0x5c7c32d83140 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d82f60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d85db0 .functor NAND 1, L_0x5c7c3312de70, L_0x5c7c3312de70, C4<1>, C4<1>;
v0x5c7c32d833b0_0 .net "in_a", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d83500_0 .net "in_b", 0 0, L_0x5c7c3312de70;  alias, 1 drivers
v0x5c7c32d835c0_0 .net "out", 0 0, L_0x5c7c32d85db0;  alias, 1 drivers
S_0x5c7c32d836c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d82f60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d83de0_0 .net "in_a", 0 0, L_0x5c7c32d85db0;  alias, 1 drivers
v0x5c7c32d83e80_0 .net "out", 0 0, L_0x5c7c3312ec10;  alias, 1 drivers
S_0x5c7c32d83890 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d836c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ec10 .functor NAND 1, L_0x5c7c32d85db0, L_0x5c7c32d85db0, C4<1>, C4<1>;
v0x5c7c32d83b00_0 .net "in_a", 0 0, L_0x5c7c32d85db0;  alias, 1 drivers
v0x5c7c32d83bf0_0 .net "in_b", 0 0, L_0x5c7c32d85db0;  alias, 1 drivers
v0x5c7c32d83ce0_0 .net "out", 0 0, L_0x5c7c3312ec10;  alias, 1 drivers
S_0x5c7c32d84380 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d81940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d853c0_0 .net "in_a", 0 0, L_0x5c7c3312ea30;  alias, 1 drivers
v0x5c7c32d85490_0 .net "in_b", 0 0, L_0x5c7c3312ecc0;  alias, 1 drivers
v0x5c7c32d85560_0 .net "out", 0 0, L_0x5c7c3312eea0;  alias, 1 drivers
v0x5c7c32d85680_0 .net "temp_out", 0 0, L_0x5c7c32d86720;  1 drivers
S_0x5c7c32d84560 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d84380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d86720 .functor NAND 1, L_0x5c7c3312ea30, L_0x5c7c3312ecc0, C4<1>, C4<1>;
v0x5c7c32d847b0_0 .net "in_a", 0 0, L_0x5c7c3312ea30;  alias, 1 drivers
v0x5c7c32d84890_0 .net "in_b", 0 0, L_0x5c7c3312ecc0;  alias, 1 drivers
v0x5c7c32d84950_0 .net "out", 0 0, L_0x5c7c32d86720;  alias, 1 drivers
S_0x5c7c32d84aa0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d84380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d85210_0 .net "in_a", 0 0, L_0x5c7c32d86720;  alias, 1 drivers
v0x5c7c32d852b0_0 .net "out", 0 0, L_0x5c7c3312eea0;  alias, 1 drivers
S_0x5c7c32d84cc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d84aa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312eea0 .functor NAND 1, L_0x5c7c32d86720, L_0x5c7c32d86720, C4<1>, C4<1>;
v0x5c7c32d84f30_0 .net "in_a", 0 0, L_0x5c7c32d86720;  alias, 1 drivers
v0x5c7c32d85020_0 .net "in_b", 0 0, L_0x5c7c32d86720;  alias, 1 drivers
v0x5c7c32d85110_0 .net "out", 0 0, L_0x5c7c3312eea0;  alias, 1 drivers
S_0x5c7c32d857d0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d81940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d85f00_0 .net "in_a", 0 0, L_0x5c7c3312e980;  alias, 1 drivers
v0x5c7c32d85fa0_0 .net "out", 0 0, L_0x5c7c3312ea30;  alias, 1 drivers
S_0x5c7c32d859a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d857d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ea30 .functor NAND 1, L_0x5c7c3312e980, L_0x5c7c3312e980, C4<1>, C4<1>;
v0x5c7c32d85c10_0 .net "in_a", 0 0, L_0x5c7c3312e980;  alias, 1 drivers
v0x5c7c32d85cd0_0 .net "in_b", 0 0, L_0x5c7c3312e980;  alias, 1 drivers
v0x5c7c32d85e20_0 .net "out", 0 0, L_0x5c7c3312ea30;  alias, 1 drivers
S_0x5c7c32d860a0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d81940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d86870_0 .net "in_a", 0 0, L_0x5c7c3312ec10;  alias, 1 drivers
v0x5c7c32d86910_0 .net "out", 0 0, L_0x5c7c3312ecc0;  alias, 1 drivers
S_0x5c7c32d86310 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d860a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ecc0 .functor NAND 1, L_0x5c7c3312ec10, L_0x5c7c3312ec10, C4<1>, C4<1>;
v0x5c7c32d86580_0 .net "in_a", 0 0, L_0x5c7c3312ec10;  alias, 1 drivers
v0x5c7c32d86640_0 .net "in_b", 0 0, L_0x5c7c3312ec10;  alias, 1 drivers
v0x5c7c32d86790_0 .net "out", 0 0, L_0x5c7c3312ecc0;  alias, 1 drivers
S_0x5c7c32d86a10 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d81940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d871b0_0 .net "in_a", 0 0, L_0x5c7c3312eea0;  alias, 1 drivers
v0x5c7c32d87250_0 .net "out", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
S_0x5c7c32d86c30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d86a10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312ef50 .functor NAND 1, L_0x5c7c3312eea0, L_0x5c7c3312eea0, C4<1>, C4<1>;
v0x5c7c32d86ea0_0 .net "in_a", 0 0, L_0x5c7c3312eea0;  alias, 1 drivers
v0x5c7c32d86f60_0 .net "in_b", 0 0, L_0x5c7c3312eea0;  alias, 1 drivers
v0x5c7c32d870b0_0 .net "out", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
S_0x5c7c32d88180 .scope module, "fa_gate14" "FullAdder" 2 19, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32da6550_0 .net "a", 0 0, L_0x5c7c33131720;  1 drivers
v0x5c7c32da65f0_0 .net "b", 0 0, L_0x5c7c331317c0;  1 drivers
v0x5c7c32da66b0_0 .net "c", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32da6750_0 .net "carry", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32da67f0_0 .net "sum", 0 0, L_0x5c7c33130dd0;  1 drivers
v0x5c7c32da6890_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c3312f350;  1 drivers
v0x5c7c32da6930_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c331304a0;  1 drivers
v0x5c7c32da69d0_0 .net "tmp_sum_out", 0 0, L_0x5c7c3312fea0;  1 drivers
S_0x5c7c32d883b0 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32d88180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d93f00_0 .net "a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d940b0_0 .net "b", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d94280_0 .net "carry", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32d94320_0 .net "sum", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
S_0x5c7c32d88620 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d883b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d896e0_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d897b0_0 .net "in_b", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d89880_0 .net "out", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32d899a0_0 .net "temp_out", 0 0, L_0x5c7c32d87040;  1 drivers
S_0x5c7c32d88890 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d88620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d87040 .functor NAND 1, L_0x5c7c33131720, L_0x5c7c331317c0, C4<1>, C4<1>;
v0x5c7c32d88b00_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d88be0_0 .net "in_b", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d88ca0_0 .net "out", 0 0, L_0x5c7c32d87040;  alias, 1 drivers
S_0x5c7c32d88dc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d88620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d89530_0 .net "in_a", 0 0, L_0x5c7c32d87040;  alias, 1 drivers
v0x5c7c32d895d0_0 .net "out", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
S_0x5c7c32d88fe0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d88dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f350 .functor NAND 1, L_0x5c7c32d87040, L_0x5c7c32d87040, C4<1>, C4<1>;
v0x5c7c32d89250_0 .net "in_a", 0 0, L_0x5c7c32d87040;  alias, 1 drivers
v0x5c7c32d89340_0 .net "in_b", 0 0, L_0x5c7c32d87040;  alias, 1 drivers
v0x5c7c32d89430_0 .net "out", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
S_0x5c7c32d89a60 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d883b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d93820_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d938c0_0 .net "in_b", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d93980_0 .net "out", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d93a20_0 .net "temp_a_and_out", 0 0, L_0x5c7c3312f560;  1 drivers
v0x5c7c32d93bd0_0 .net "temp_a_out", 0 0, L_0x5c7c3312f400;  1 drivers
v0x5c7c32d93c70_0 .net "temp_b_and_out", 0 0, L_0x5c7c3312f770;  1 drivers
v0x5c7c32d93e20_0 .net "temp_b_out", 0 0, L_0x5c7c3312f610;  1 drivers
S_0x5c7c32d89c40 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d89a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d8ad00_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d8ada0_0 .net "in_b", 0 0, L_0x5c7c3312f400;  alias, 1 drivers
v0x5c7c32d8ae90_0 .net "out", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
v0x5c7c32d8afb0_0 .net "temp_out", 0 0, L_0x5c7c3312f4b0;  1 drivers
S_0x5c7c32d89eb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d89c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f4b0 .functor NAND 1, L_0x5c7c33131720, L_0x5c7c3312f400, C4<1>, C4<1>;
v0x5c7c32d8a120_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d8a230_0 .net "in_b", 0 0, L_0x5c7c3312f400;  alias, 1 drivers
v0x5c7c32d8a2f0_0 .net "out", 0 0, L_0x5c7c3312f4b0;  alias, 1 drivers
S_0x5c7c32d8a410 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d89c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d8ab50_0 .net "in_a", 0 0, L_0x5c7c3312f4b0;  alias, 1 drivers
v0x5c7c32d8abf0_0 .net "out", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
S_0x5c7c32d8a630 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d8a410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f560 .functor NAND 1, L_0x5c7c3312f4b0, L_0x5c7c3312f4b0, C4<1>, C4<1>;
v0x5c7c32d8a8a0_0 .net "in_a", 0 0, L_0x5c7c3312f4b0;  alias, 1 drivers
v0x5c7c32d8a960_0 .net "in_b", 0 0, L_0x5c7c3312f4b0;  alias, 1 drivers
v0x5c7c32d8aa50_0 .net "out", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
S_0x5c7c32d8b070 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d89a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d8c0a0_0 .net "in_a", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d8c140_0 .net "in_b", 0 0, L_0x5c7c3312f610;  alias, 1 drivers
v0x5c7c32d8c230_0 .net "out", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
v0x5c7c32d8c350_0 .net "temp_out", 0 0, L_0x5c7c3312f6c0;  1 drivers
S_0x5c7c32d8b250 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d8b070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f6c0 .functor NAND 1, L_0x5c7c331317c0, L_0x5c7c3312f610, C4<1>, C4<1>;
v0x5c7c32d8b4c0_0 .net "in_a", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d8b5d0_0 .net "in_b", 0 0, L_0x5c7c3312f610;  alias, 1 drivers
v0x5c7c32d8b690_0 .net "out", 0 0, L_0x5c7c3312f6c0;  alias, 1 drivers
S_0x5c7c32d8b7b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d8b070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d8bef0_0 .net "in_a", 0 0, L_0x5c7c3312f6c0;  alias, 1 drivers
v0x5c7c32d8bf90_0 .net "out", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
S_0x5c7c32d8b9d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d8b7b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f770 .functor NAND 1, L_0x5c7c3312f6c0, L_0x5c7c3312f6c0, C4<1>, C4<1>;
v0x5c7c32d8bc40_0 .net "in_a", 0 0, L_0x5c7c3312f6c0;  alias, 1 drivers
v0x5c7c32d8bd00_0 .net "in_b", 0 0, L_0x5c7c3312f6c0;  alias, 1 drivers
v0x5c7c32d8bdf0_0 .net "out", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
S_0x5c7c32d8c4a0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d89a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d8cbe0_0 .net "in_a", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d8cc80_0 .net "out", 0 0, L_0x5c7c3312f400;  alias, 1 drivers
S_0x5c7c32d8c670 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d8c4a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f400 .functor NAND 1, L_0x5c7c331317c0, L_0x5c7c331317c0, C4<1>, C4<1>;
v0x5c7c32d8c8c0_0 .net "in_a", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d8ca10_0 .net "in_b", 0 0, L_0x5c7c331317c0;  alias, 1 drivers
v0x5c7c32d8cad0_0 .net "out", 0 0, L_0x5c7c3312f400;  alias, 1 drivers
S_0x5c7c32d8cd80 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d89a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d8d500_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d8d5a0_0 .net "out", 0 0, L_0x5c7c3312f610;  alias, 1 drivers
S_0x5c7c32d8cfa0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d8cd80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f610 .functor NAND 1, L_0x5c7c33131720, L_0x5c7c33131720, C4<1>, C4<1>;
v0x5c7c32d8d210_0 .net "in_a", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d8d360_0 .net "in_b", 0 0, L_0x5c7c33131720;  alias, 1 drivers
v0x5c7c32d8d420_0 .net "out", 0 0, L_0x5c7c3312f610;  alias, 1 drivers
S_0x5c7c32d8d6a0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d89a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d93170_0 .net "branch1_out", 0 0, L_0x5c7c3312f980;  1 drivers
v0x5c7c32d932a0_0 .net "branch2_out", 0 0, L_0x5c7c3312fc10;  1 drivers
v0x5c7c32d933f0_0 .net "in_a", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
v0x5c7c32d934c0_0 .net "in_b", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
v0x5c7c32d93560_0 .net "out", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d93600_0 .net "temp1_out", 0 0, L_0x5c7c3312f8d0;  1 drivers
v0x5c7c32d936a0_0 .net "temp2_out", 0 0, L_0x5c7c3312fb60;  1 drivers
v0x5c7c32d93740_0 .net "temp3_out", 0 0, L_0x5c7c3312fdf0;  1 drivers
S_0x5c7c32d8d920 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d8d6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d8e9b0_0 .net "in_a", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
v0x5c7c32d8ea50_0 .net "in_b", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
v0x5c7c32d8eb10_0 .net "out", 0 0, L_0x5c7c3312f8d0;  alias, 1 drivers
v0x5c7c32d8ec30_0 .net "temp_out", 0 0, L_0x5c7c3312f820;  1 drivers
S_0x5c7c32d8db90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d8d920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f820 .functor NAND 1, L_0x5c7c3312f560, L_0x5c7c3312f560, C4<1>, C4<1>;
v0x5c7c32d8de00_0 .net "in_a", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
v0x5c7c32d8dec0_0 .net "in_b", 0 0, L_0x5c7c3312f560;  alias, 1 drivers
v0x5c7c32d8e010_0 .net "out", 0 0, L_0x5c7c3312f820;  alias, 1 drivers
S_0x5c7c32d8e110 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d8d920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d8e800_0 .net "in_a", 0 0, L_0x5c7c3312f820;  alias, 1 drivers
v0x5c7c32d8e8a0_0 .net "out", 0 0, L_0x5c7c3312f8d0;  alias, 1 drivers
S_0x5c7c32d8e2e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d8e110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f8d0 .functor NAND 1, L_0x5c7c3312f820, L_0x5c7c3312f820, C4<1>, C4<1>;
v0x5c7c32d8e550_0 .net "in_a", 0 0, L_0x5c7c3312f820;  alias, 1 drivers
v0x5c7c32d8e610_0 .net "in_b", 0 0, L_0x5c7c3312f820;  alias, 1 drivers
v0x5c7c32d8e700_0 .net "out", 0 0, L_0x5c7c3312f8d0;  alias, 1 drivers
S_0x5c7c32d8eda0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d8d6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d8fdd0_0 .net "in_a", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
v0x5c7c32d8fe70_0 .net "in_b", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
v0x5c7c32d8ff30_0 .net "out", 0 0, L_0x5c7c3312fb60;  alias, 1 drivers
v0x5c7c32d90050_0 .net "temp_out", 0 0, L_0x5c7c32d91bf0;  1 drivers
S_0x5c7c32d8ef80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d8eda0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d91bf0 .functor NAND 1, L_0x5c7c3312f770, L_0x5c7c3312f770, C4<1>, C4<1>;
v0x5c7c32d8f1f0_0 .net "in_a", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
v0x5c7c32d8f2b0_0 .net "in_b", 0 0, L_0x5c7c3312f770;  alias, 1 drivers
v0x5c7c32d8f400_0 .net "out", 0 0, L_0x5c7c32d91bf0;  alias, 1 drivers
S_0x5c7c32d8f500 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d8eda0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d8fc20_0 .net "in_a", 0 0, L_0x5c7c32d91bf0;  alias, 1 drivers
v0x5c7c32d8fcc0_0 .net "out", 0 0, L_0x5c7c3312fb60;  alias, 1 drivers
S_0x5c7c32d8f6d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d8f500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312fb60 .functor NAND 1, L_0x5c7c32d91bf0, L_0x5c7c32d91bf0, C4<1>, C4<1>;
v0x5c7c32d8f940_0 .net "in_a", 0 0, L_0x5c7c32d91bf0;  alias, 1 drivers
v0x5c7c32d8fa30_0 .net "in_b", 0 0, L_0x5c7c32d91bf0;  alias, 1 drivers
v0x5c7c32d8fb20_0 .net "out", 0 0, L_0x5c7c3312fb60;  alias, 1 drivers
S_0x5c7c32d901c0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d8d6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d91200_0 .net "in_a", 0 0, L_0x5c7c3312f980;  alias, 1 drivers
v0x5c7c32d912d0_0 .net "in_b", 0 0, L_0x5c7c3312fc10;  alias, 1 drivers
v0x5c7c32d913a0_0 .net "out", 0 0, L_0x5c7c3312fdf0;  alias, 1 drivers
v0x5c7c32d914c0_0 .net "temp_out", 0 0, L_0x5c7c32d92560;  1 drivers
S_0x5c7c32d903a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d901c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d92560 .functor NAND 1, L_0x5c7c3312f980, L_0x5c7c3312fc10, C4<1>, C4<1>;
v0x5c7c32d905f0_0 .net "in_a", 0 0, L_0x5c7c3312f980;  alias, 1 drivers
v0x5c7c32d906d0_0 .net "in_b", 0 0, L_0x5c7c3312fc10;  alias, 1 drivers
v0x5c7c32d90790_0 .net "out", 0 0, L_0x5c7c32d92560;  alias, 1 drivers
S_0x5c7c32d908e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d901c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d91050_0 .net "in_a", 0 0, L_0x5c7c32d92560;  alias, 1 drivers
v0x5c7c32d910f0_0 .net "out", 0 0, L_0x5c7c3312fdf0;  alias, 1 drivers
S_0x5c7c32d90b00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d908e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312fdf0 .functor NAND 1, L_0x5c7c32d92560, L_0x5c7c32d92560, C4<1>, C4<1>;
v0x5c7c32d90d70_0 .net "in_a", 0 0, L_0x5c7c32d92560;  alias, 1 drivers
v0x5c7c32d90e60_0 .net "in_b", 0 0, L_0x5c7c32d92560;  alias, 1 drivers
v0x5c7c32d90f50_0 .net "out", 0 0, L_0x5c7c3312fdf0;  alias, 1 drivers
S_0x5c7c32d91610 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d8d6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d91d40_0 .net "in_a", 0 0, L_0x5c7c3312f8d0;  alias, 1 drivers
v0x5c7c32d91de0_0 .net "out", 0 0, L_0x5c7c3312f980;  alias, 1 drivers
S_0x5c7c32d917e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d91610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312f980 .functor NAND 1, L_0x5c7c3312f8d0, L_0x5c7c3312f8d0, C4<1>, C4<1>;
v0x5c7c32d91a50_0 .net "in_a", 0 0, L_0x5c7c3312f8d0;  alias, 1 drivers
v0x5c7c32d91b10_0 .net "in_b", 0 0, L_0x5c7c3312f8d0;  alias, 1 drivers
v0x5c7c32d91c60_0 .net "out", 0 0, L_0x5c7c3312f980;  alias, 1 drivers
S_0x5c7c32d91ee0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d8d6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d926b0_0 .net "in_a", 0 0, L_0x5c7c3312fb60;  alias, 1 drivers
v0x5c7c32d92750_0 .net "out", 0 0, L_0x5c7c3312fc10;  alias, 1 drivers
S_0x5c7c32d92150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d91ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312fc10 .functor NAND 1, L_0x5c7c3312fb60, L_0x5c7c3312fb60, C4<1>, C4<1>;
v0x5c7c32d923c0_0 .net "in_a", 0 0, L_0x5c7c3312fb60;  alias, 1 drivers
v0x5c7c32d92480_0 .net "in_b", 0 0, L_0x5c7c3312fb60;  alias, 1 drivers
v0x5c7c32d925d0_0 .net "out", 0 0, L_0x5c7c3312fc10;  alias, 1 drivers
S_0x5c7c32d92850 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d8d6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d92ff0_0 .net "in_a", 0 0, L_0x5c7c3312fdf0;  alias, 1 drivers
v0x5c7c32d93090_0 .net "out", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
S_0x5c7c32d92a70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d92850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3312fea0 .functor NAND 1, L_0x5c7c3312fdf0, L_0x5c7c3312fdf0, C4<1>, C4<1>;
v0x5c7c32d92ce0_0 .net "in_a", 0 0, L_0x5c7c3312fdf0;  alias, 1 drivers
v0x5c7c32d92da0_0 .net "in_b", 0 0, L_0x5c7c3312fdf0;  alias, 1 drivers
v0x5c7c32d92ef0_0 .net "out", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
S_0x5c7c32d94400 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32d88180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32d9ff20_0 .net "a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d9ffc0_0 .net "b", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32da0080_0 .net "carry", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32da0120_0 .net "sum", 0 0, L_0x5c7c33130dd0;  alias, 1 drivers
S_0x5c7c32d94620 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32d94400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d955c0_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d95660_0 .net "in_b", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d95720_0 .net "out", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32d95840_0 .net "temp_out", 0 0, L_0x5c7c32d92e80;  1 drivers
S_0x5c7c32d947d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d94620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d92e80 .functor NAND 1, L_0x5c7c3312fea0, L_0x5c7c3312ef50, C4<1>, C4<1>;
v0x5c7c32d94a40_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d94b00_0 .net "in_b", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d94bc0_0 .net "out", 0 0, L_0x5c7c32d92e80;  alias, 1 drivers
S_0x5c7c32d94cf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d94620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d95410_0 .net "in_a", 0 0, L_0x5c7c32d92e80;  alias, 1 drivers
v0x5c7c32d954b0_0 .net "out", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
S_0x5c7c32d94ec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d94cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331304a0 .functor NAND 1, L_0x5c7c32d92e80, L_0x5c7c32d92e80, C4<1>, C4<1>;
v0x5c7c32d95130_0 .net "in_a", 0 0, L_0x5c7c32d92e80;  alias, 1 drivers
v0x5c7c32d95220_0 .net "in_b", 0 0, L_0x5c7c32d92e80;  alias, 1 drivers
v0x5c7c32d95310_0 .net "out", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
S_0x5c7c32d959b0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32d94400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d9f840_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d9f8e0_0 .net "in_b", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d9f9a0_0 .net "out", 0 0, L_0x5c7c33130dd0;  alias, 1 drivers
v0x5c7c32d9fa40_0 .net "temp_a_and_out", 0 0, L_0x5c7c331306b0;  1 drivers
v0x5c7c32d9fbf0_0 .net "temp_a_out", 0 0, L_0x5c7c33130550;  1 drivers
v0x5c7c32d9fc90_0 .net "temp_b_and_out", 0 0, L_0x5c7c331308c0;  1 drivers
v0x5c7c32d9fe40_0 .net "temp_b_out", 0 0, L_0x5c7c33130760;  1 drivers
S_0x5c7c32d95b90 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32d959b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d96c30_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d96de0_0 .net "in_b", 0 0, L_0x5c7c33130550;  alias, 1 drivers
v0x5c7c32d96ed0_0 .net "out", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
v0x5c7c32d96ff0_0 .net "temp_out", 0 0, L_0x5c7c33130600;  1 drivers
S_0x5c7c32d95e00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d95b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130600 .functor NAND 1, L_0x5c7c3312fea0, L_0x5c7c33130550, C4<1>, C4<1>;
v0x5c7c32d96070_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d96130_0 .net "in_b", 0 0, L_0x5c7c33130550;  alias, 1 drivers
v0x5c7c32d961f0_0 .net "out", 0 0, L_0x5c7c33130600;  alias, 1 drivers
S_0x5c7c32d96310 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d95b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d96a80_0 .net "in_a", 0 0, L_0x5c7c33130600;  alias, 1 drivers
v0x5c7c32d96b20_0 .net "out", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
S_0x5c7c32d96530 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d96310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331306b0 .functor NAND 1, L_0x5c7c33130600, L_0x5c7c33130600, C4<1>, C4<1>;
v0x5c7c32d967a0_0 .net "in_a", 0 0, L_0x5c7c33130600;  alias, 1 drivers
v0x5c7c32d96890_0 .net "in_b", 0 0, L_0x5c7c33130600;  alias, 1 drivers
v0x5c7c32d96980_0 .net "out", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
S_0x5c7c32d970b0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32d959b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d980c0_0 .net "in_a", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d98160_0 .net "in_b", 0 0, L_0x5c7c33130760;  alias, 1 drivers
v0x5c7c32d98250_0 .net "out", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
v0x5c7c32d98370_0 .net "temp_out", 0 0, L_0x5c7c33130810;  1 drivers
S_0x5c7c32d97290 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d970b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130810 .functor NAND 1, L_0x5c7c3312ef50, L_0x5c7c33130760, C4<1>, C4<1>;
v0x5c7c32d97500_0 .net "in_a", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d975c0_0 .net "in_b", 0 0, L_0x5c7c33130760;  alias, 1 drivers
v0x5c7c32d97680_0 .net "out", 0 0, L_0x5c7c33130810;  alias, 1 drivers
S_0x5c7c32d977a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d970b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d97f10_0 .net "in_a", 0 0, L_0x5c7c33130810;  alias, 1 drivers
v0x5c7c32d97fb0_0 .net "out", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
S_0x5c7c32d979c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d977a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331308c0 .functor NAND 1, L_0x5c7c33130810, L_0x5c7c33130810, C4<1>, C4<1>;
v0x5c7c32d97c30_0 .net "in_a", 0 0, L_0x5c7c33130810;  alias, 1 drivers
v0x5c7c32d97d20_0 .net "in_b", 0 0, L_0x5c7c33130810;  alias, 1 drivers
v0x5c7c32d97e10_0 .net "out", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
S_0x5c7c32d984c0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32d959b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d98cd0_0 .net "in_a", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d98d70_0 .net "out", 0 0, L_0x5c7c33130550;  alias, 1 drivers
S_0x5c7c32d98690 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d984c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130550 .functor NAND 1, L_0x5c7c3312ef50, L_0x5c7c3312ef50, C4<1>, C4<1>;
v0x5c7c32d988e0_0 .net "in_a", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d98ab0_0 .net "in_b", 0 0, L_0x5c7c3312ef50;  alias, 1 drivers
v0x5c7c32d98b70_0 .net "out", 0 0, L_0x5c7c33130550;  alias, 1 drivers
S_0x5c7c32d98e70 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32d959b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d995b0_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d99650_0 .net "out", 0 0, L_0x5c7c33130760;  alias, 1 drivers
S_0x5c7c32d99090 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d98e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130760 .functor NAND 1, L_0x5c7c3312fea0, L_0x5c7c3312fea0, C4<1>, C4<1>;
v0x5c7c32d99300_0 .net "in_a", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d993c0_0 .net "in_b", 0 0, L_0x5c7c3312fea0;  alias, 1 drivers
v0x5c7c32d99480_0 .net "out", 0 0, L_0x5c7c33130760;  alias, 1 drivers
S_0x5c7c32d99750 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32d959b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d9f190_0 .net "branch1_out", 0 0, L_0x5c7c33130ad0;  1 drivers
v0x5c7c32d9f2c0_0 .net "branch2_out", 0 0, L_0x5c7c33130c50;  1 drivers
v0x5c7c32d9f410_0 .net "in_a", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
v0x5c7c32d9f4e0_0 .net "in_b", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
v0x5c7c32d9f580_0 .net "out", 0 0, L_0x5c7c33130dd0;  alias, 1 drivers
v0x5c7c32d9f620_0 .net "temp1_out", 0 0, L_0x5c7c33130a20;  1 drivers
v0x5c7c32d9f6c0_0 .net "temp2_out", 0 0, L_0x5c7c33130ba0;  1 drivers
v0x5c7c32d9f760_0 .net "temp3_out", 0 0, L_0x5c7c33130d20;  1 drivers
S_0x5c7c32d999d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32d99750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d9a9d0_0 .net "in_a", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
v0x5c7c32d9aa70_0 .net "in_b", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
v0x5c7c32d9ab30_0 .net "out", 0 0, L_0x5c7c33130a20;  alias, 1 drivers
v0x5c7c32d9ac50_0 .net "temp_out", 0 0, L_0x5c7c33130970;  1 drivers
S_0x5c7c32d99c40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d999d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130970 .functor NAND 1, L_0x5c7c331306b0, L_0x5c7c331306b0, C4<1>, C4<1>;
v0x5c7c32d99eb0_0 .net "in_a", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
v0x5c7c32d99f70_0 .net "in_b", 0 0, L_0x5c7c331306b0;  alias, 1 drivers
v0x5c7c32d9a030_0 .net "out", 0 0, L_0x5c7c33130970;  alias, 1 drivers
S_0x5c7c32d9a130 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d999d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d9a820_0 .net "in_a", 0 0, L_0x5c7c33130970;  alias, 1 drivers
v0x5c7c32d9a8c0_0 .net "out", 0 0, L_0x5c7c33130a20;  alias, 1 drivers
S_0x5c7c32d9a300 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d9a130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130a20 .functor NAND 1, L_0x5c7c33130970, L_0x5c7c33130970, C4<1>, C4<1>;
v0x5c7c32d9a570_0 .net "in_a", 0 0, L_0x5c7c33130970;  alias, 1 drivers
v0x5c7c32d9a630_0 .net "in_b", 0 0, L_0x5c7c33130970;  alias, 1 drivers
v0x5c7c32d9a720_0 .net "out", 0 0, L_0x5c7c33130a20;  alias, 1 drivers
S_0x5c7c32d9adc0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32d99750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d9bdf0_0 .net "in_a", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
v0x5c7c32d9be90_0 .net "in_b", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
v0x5c7c32d9bf50_0 .net "out", 0 0, L_0x5c7c33130ba0;  alias, 1 drivers
v0x5c7c32d9c070_0 .net "temp_out", 0 0, L_0x5c7c32d9dc10;  1 drivers
S_0x5c7c32d9afa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d9adc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d9dc10 .functor NAND 1, L_0x5c7c331308c0, L_0x5c7c331308c0, C4<1>, C4<1>;
v0x5c7c32d9b210_0 .net "in_a", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
v0x5c7c32d9b2d0_0 .net "in_b", 0 0, L_0x5c7c331308c0;  alias, 1 drivers
v0x5c7c32d9b420_0 .net "out", 0 0, L_0x5c7c32d9dc10;  alias, 1 drivers
S_0x5c7c32d9b520 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d9adc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d9bc40_0 .net "in_a", 0 0, L_0x5c7c32d9dc10;  alias, 1 drivers
v0x5c7c32d9bce0_0 .net "out", 0 0, L_0x5c7c33130ba0;  alias, 1 drivers
S_0x5c7c32d9b6f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d9b520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130ba0 .functor NAND 1, L_0x5c7c32d9dc10, L_0x5c7c32d9dc10, C4<1>, C4<1>;
v0x5c7c32d9b960_0 .net "in_a", 0 0, L_0x5c7c32d9dc10;  alias, 1 drivers
v0x5c7c32d9ba50_0 .net "in_b", 0 0, L_0x5c7c32d9dc10;  alias, 1 drivers
v0x5c7c32d9bb40_0 .net "out", 0 0, L_0x5c7c33130ba0;  alias, 1 drivers
S_0x5c7c32d9c1e0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32d99750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32d9d220_0 .net "in_a", 0 0, L_0x5c7c33130ad0;  alias, 1 drivers
v0x5c7c32d9d2f0_0 .net "in_b", 0 0, L_0x5c7c33130c50;  alias, 1 drivers
v0x5c7c32d9d3c0_0 .net "out", 0 0, L_0x5c7c33130d20;  alias, 1 drivers
v0x5c7c32d9d4e0_0 .net "temp_out", 0 0, L_0x5c7c32d9e580;  1 drivers
S_0x5c7c32d9c3c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32d9c1e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d9e580 .functor NAND 1, L_0x5c7c33130ad0, L_0x5c7c33130c50, C4<1>, C4<1>;
v0x5c7c32d9c610_0 .net "in_a", 0 0, L_0x5c7c33130ad0;  alias, 1 drivers
v0x5c7c32d9c6f0_0 .net "in_b", 0 0, L_0x5c7c33130c50;  alias, 1 drivers
v0x5c7c32d9c7b0_0 .net "out", 0 0, L_0x5c7c32d9e580;  alias, 1 drivers
S_0x5c7c32d9c900 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32d9c1e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d9d070_0 .net "in_a", 0 0, L_0x5c7c32d9e580;  alias, 1 drivers
v0x5c7c32d9d110_0 .net "out", 0 0, L_0x5c7c33130d20;  alias, 1 drivers
S_0x5c7c32d9cb20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d9c900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130d20 .functor NAND 1, L_0x5c7c32d9e580, L_0x5c7c32d9e580, C4<1>, C4<1>;
v0x5c7c32d9cd90_0 .net "in_a", 0 0, L_0x5c7c32d9e580;  alias, 1 drivers
v0x5c7c32d9ce80_0 .net "in_b", 0 0, L_0x5c7c32d9e580;  alias, 1 drivers
v0x5c7c32d9cf70_0 .net "out", 0 0, L_0x5c7c33130d20;  alias, 1 drivers
S_0x5c7c32d9d630 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32d99750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d9dd60_0 .net "in_a", 0 0, L_0x5c7c33130a20;  alias, 1 drivers
v0x5c7c32d9de00_0 .net "out", 0 0, L_0x5c7c33130ad0;  alias, 1 drivers
S_0x5c7c32d9d800 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d9d630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130ad0 .functor NAND 1, L_0x5c7c33130a20, L_0x5c7c33130a20, C4<1>, C4<1>;
v0x5c7c32d9da70_0 .net "in_a", 0 0, L_0x5c7c33130a20;  alias, 1 drivers
v0x5c7c32d9db30_0 .net "in_b", 0 0, L_0x5c7c33130a20;  alias, 1 drivers
v0x5c7c32d9dc80_0 .net "out", 0 0, L_0x5c7c33130ad0;  alias, 1 drivers
S_0x5c7c32d9df00 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32d99750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d9e6d0_0 .net "in_a", 0 0, L_0x5c7c33130ba0;  alias, 1 drivers
v0x5c7c32d9e770_0 .net "out", 0 0, L_0x5c7c33130c50;  alias, 1 drivers
S_0x5c7c32d9e170 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d9df00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130c50 .functor NAND 1, L_0x5c7c33130ba0, L_0x5c7c33130ba0, C4<1>, C4<1>;
v0x5c7c32d9e3e0_0 .net "in_a", 0 0, L_0x5c7c33130ba0;  alias, 1 drivers
v0x5c7c32d9e4a0_0 .net "in_b", 0 0, L_0x5c7c33130ba0;  alias, 1 drivers
v0x5c7c32d9e5f0_0 .net "out", 0 0, L_0x5c7c33130c50;  alias, 1 drivers
S_0x5c7c32d9e870 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32d99750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32d9f010_0 .net "in_a", 0 0, L_0x5c7c33130d20;  alias, 1 drivers
v0x5c7c32d9f0b0_0 .net "out", 0 0, L_0x5c7c33130dd0;  alias, 1 drivers
S_0x5c7c32d9ea90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32d9e870;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130dd0 .functor NAND 1, L_0x5c7c33130d20, L_0x5c7c33130d20, C4<1>, C4<1>;
v0x5c7c32d9ed00_0 .net "in_a", 0 0, L_0x5c7c33130d20;  alias, 1 drivers
v0x5c7c32d9edc0_0 .net "in_b", 0 0, L_0x5c7c33130d20;  alias, 1 drivers
v0x5c7c32d9ef10_0 .net "out", 0 0, L_0x5c7c33130dd0;  alias, 1 drivers
S_0x5c7c32da0290 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32d88180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32da5c80_0 .net "branch1_out", 0 0, L_0x5c7c33131060;  1 drivers
v0x5c7c32da5db0_0 .net "branch2_out", 0 0, L_0x5c7c331312f0;  1 drivers
v0x5c7c32da5f00_0 .net "in_a", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32da60e0_0 .net "in_b", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32da6290_0 .net "out", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32da6330_0 .net "temp1_out", 0 0, L_0x5c7c33130fb0;  1 drivers
v0x5c7c32da63d0_0 .net "temp2_out", 0 0, L_0x5c7c33131240;  1 drivers
v0x5c7c32da6470_0 .net "temp3_out", 0 0, L_0x5c7c331314d0;  1 drivers
S_0x5c7c32da0420 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32da0290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32da14c0_0 .net "in_a", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32da1560_0 .net "in_b", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32da1620_0 .net "out", 0 0, L_0x5c7c33130fb0;  alias, 1 drivers
v0x5c7c32da1740_0 .net "temp_out", 0 0, L_0x5c7c32d9eea0;  1 drivers
S_0x5c7c32da0640 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32da0420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32d9eea0 .functor NAND 1, L_0x5c7c3312f350, L_0x5c7c3312f350, C4<1>, C4<1>;
v0x5c7c32da08b0_0 .net "in_a", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32da0a00_0 .net "in_b", 0 0, L_0x5c7c3312f350;  alias, 1 drivers
v0x5c7c32da0ac0_0 .net "out", 0 0, L_0x5c7c32d9eea0;  alias, 1 drivers
S_0x5c7c32da0bf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32da0420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da1310_0 .net "in_a", 0 0, L_0x5c7c32d9eea0;  alias, 1 drivers
v0x5c7c32da13b0_0 .net "out", 0 0, L_0x5c7c33130fb0;  alias, 1 drivers
S_0x5c7c32da0dc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da0bf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33130fb0 .functor NAND 1, L_0x5c7c32d9eea0, L_0x5c7c32d9eea0, C4<1>, C4<1>;
v0x5c7c32da1030_0 .net "in_a", 0 0, L_0x5c7c32d9eea0;  alias, 1 drivers
v0x5c7c32da1120_0 .net "in_b", 0 0, L_0x5c7c32d9eea0;  alias, 1 drivers
v0x5c7c32da1210_0 .net "out", 0 0, L_0x5c7c33130fb0;  alias, 1 drivers
S_0x5c7c32da18b0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32da0290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32da28e0_0 .net "in_a", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32da2980_0 .net "in_b", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32da2a40_0 .net "out", 0 0, L_0x5c7c33131240;  alias, 1 drivers
v0x5c7c32da2b60_0 .net "temp_out", 0 0, L_0x5c7c32da4700;  1 drivers
S_0x5c7c32da1a90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32da18b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32da4700 .functor NAND 1, L_0x5c7c331304a0, L_0x5c7c331304a0, C4<1>, C4<1>;
v0x5c7c32da1d00_0 .net "in_a", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32da1e50_0 .net "in_b", 0 0, L_0x5c7c331304a0;  alias, 1 drivers
v0x5c7c32da1f10_0 .net "out", 0 0, L_0x5c7c32da4700;  alias, 1 drivers
S_0x5c7c32da2010 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32da18b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da2730_0 .net "in_a", 0 0, L_0x5c7c32da4700;  alias, 1 drivers
v0x5c7c32da27d0_0 .net "out", 0 0, L_0x5c7c33131240;  alias, 1 drivers
S_0x5c7c32da21e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da2010;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131240 .functor NAND 1, L_0x5c7c32da4700, L_0x5c7c32da4700, C4<1>, C4<1>;
v0x5c7c32da2450_0 .net "in_a", 0 0, L_0x5c7c32da4700;  alias, 1 drivers
v0x5c7c32da2540_0 .net "in_b", 0 0, L_0x5c7c32da4700;  alias, 1 drivers
v0x5c7c32da2630_0 .net "out", 0 0, L_0x5c7c33131240;  alias, 1 drivers
S_0x5c7c32da2cd0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32da0290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32da3d10_0 .net "in_a", 0 0, L_0x5c7c33131060;  alias, 1 drivers
v0x5c7c32da3de0_0 .net "in_b", 0 0, L_0x5c7c331312f0;  alias, 1 drivers
v0x5c7c32da3eb0_0 .net "out", 0 0, L_0x5c7c331314d0;  alias, 1 drivers
v0x5c7c32da3fd0_0 .net "temp_out", 0 0, L_0x5c7c32da5070;  1 drivers
S_0x5c7c32da2eb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32da2cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32da5070 .functor NAND 1, L_0x5c7c33131060, L_0x5c7c331312f0, C4<1>, C4<1>;
v0x5c7c32da3100_0 .net "in_a", 0 0, L_0x5c7c33131060;  alias, 1 drivers
v0x5c7c32da31e0_0 .net "in_b", 0 0, L_0x5c7c331312f0;  alias, 1 drivers
v0x5c7c32da32a0_0 .net "out", 0 0, L_0x5c7c32da5070;  alias, 1 drivers
S_0x5c7c32da33f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32da2cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da3b60_0 .net "in_a", 0 0, L_0x5c7c32da5070;  alias, 1 drivers
v0x5c7c32da3c00_0 .net "out", 0 0, L_0x5c7c331314d0;  alias, 1 drivers
S_0x5c7c32da3610 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da33f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331314d0 .functor NAND 1, L_0x5c7c32da5070, L_0x5c7c32da5070, C4<1>, C4<1>;
v0x5c7c32da3880_0 .net "in_a", 0 0, L_0x5c7c32da5070;  alias, 1 drivers
v0x5c7c32da3970_0 .net "in_b", 0 0, L_0x5c7c32da5070;  alias, 1 drivers
v0x5c7c32da3a60_0 .net "out", 0 0, L_0x5c7c331314d0;  alias, 1 drivers
S_0x5c7c32da4120 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32da0290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da4850_0 .net "in_a", 0 0, L_0x5c7c33130fb0;  alias, 1 drivers
v0x5c7c32da48f0_0 .net "out", 0 0, L_0x5c7c33131060;  alias, 1 drivers
S_0x5c7c32da42f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da4120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131060 .functor NAND 1, L_0x5c7c33130fb0, L_0x5c7c33130fb0, C4<1>, C4<1>;
v0x5c7c32da4560_0 .net "in_a", 0 0, L_0x5c7c33130fb0;  alias, 1 drivers
v0x5c7c32da4620_0 .net "in_b", 0 0, L_0x5c7c33130fb0;  alias, 1 drivers
v0x5c7c32da4770_0 .net "out", 0 0, L_0x5c7c33131060;  alias, 1 drivers
S_0x5c7c32da49f0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32da0290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da51c0_0 .net "in_a", 0 0, L_0x5c7c33131240;  alias, 1 drivers
v0x5c7c32da5260_0 .net "out", 0 0, L_0x5c7c331312f0;  alias, 1 drivers
S_0x5c7c32da4c60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da49f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331312f0 .functor NAND 1, L_0x5c7c33131240, L_0x5c7c33131240, C4<1>, C4<1>;
v0x5c7c32da4ed0_0 .net "in_a", 0 0, L_0x5c7c33131240;  alias, 1 drivers
v0x5c7c32da4f90_0 .net "in_b", 0 0, L_0x5c7c33131240;  alias, 1 drivers
v0x5c7c32da50e0_0 .net "out", 0 0, L_0x5c7c331312f0;  alias, 1 drivers
S_0x5c7c32da5360 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32da0290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da5b00_0 .net "in_a", 0 0, L_0x5c7c331314d0;  alias, 1 drivers
v0x5c7c32da5ba0_0 .net "out", 0 0, L_0x5c7c33131580;  alias, 1 drivers
S_0x5c7c32da5580 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da5360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131580 .functor NAND 1, L_0x5c7c331314d0, L_0x5c7c331314d0, C4<1>, C4<1>;
v0x5c7c32da57f0_0 .net "in_a", 0 0, L_0x5c7c331314d0;  alias, 1 drivers
v0x5c7c32da58b0_0 .net "in_b", 0 0, L_0x5c7c331314d0;  alias, 1 drivers
v0x5c7c32da5a00_0 .net "out", 0 0, L_0x5c7c33131580;  alias, 1 drivers
S_0x5c7c32da6ad0 .scope module, "fa_gate15" "FullAdder" 2 20, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32dc4e80_0 .net "a", 0 0, L_0x5c7c33133d60;  1 drivers
v0x5c7c32dc4f20_0 .net "b", 0 0, L_0x5c7c33133e00;  1 drivers
v0x5c7c32dc4fe0_0 .net "c", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32dc5080_0 .net "carry", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dc5120_0 .net "sum", 0 0, L_0x5c7c33133410;  1 drivers
v0x5c7c32dc51c0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33131990;  1 drivers
v0x5c7c32dc5260_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33132ae0;  1 drivers
v0x5c7c32dc5300_0 .net "tmp_sum_out", 0 0, L_0x5c7c331324e0;  1 drivers
S_0x5c7c32da6cb0 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32da6ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32db2830_0 .net "a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32db29e0_0 .net "b", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32db2bb0_0 .net "carry", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32db2c50_0 .net "sum", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
S_0x5c7c32da6f20 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32da6cb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32da8010_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32da80e0_0 .net "in_b", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32da81b0_0 .net "out", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32da82d0_0 .net "temp_out", 0 0, L_0x5c7c32da5990;  1 drivers
S_0x5c7c32da7190 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32da6f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32da5990 .functor NAND 1, L_0x5c7c33133d60, L_0x5c7c33133e00, C4<1>, C4<1>;
v0x5c7c32da7400_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32da74e0_0 .net "in_b", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32da75a0_0 .net "out", 0 0, L_0x5c7c32da5990;  alias, 1 drivers
S_0x5c7c32da76f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32da6f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da7e60_0 .net "in_a", 0 0, L_0x5c7c32da5990;  alias, 1 drivers
v0x5c7c32da7f00_0 .net "out", 0 0, L_0x5c7c33131990;  alias, 1 drivers
S_0x5c7c32da7910 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da76f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131990 .functor NAND 1, L_0x5c7c32da5990, L_0x5c7c32da5990, C4<1>, C4<1>;
v0x5c7c32da7b80_0 .net "in_a", 0 0, L_0x5c7c32da5990;  alias, 1 drivers
v0x5c7c32da7c70_0 .net "in_b", 0 0, L_0x5c7c32da5990;  alias, 1 drivers
v0x5c7c32da7d60_0 .net "out", 0 0, L_0x5c7c33131990;  alias, 1 drivers
S_0x5c7c32da8390 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32da6cb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32db2150_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32db21f0_0 .net "in_b", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32db22b0_0 .net "out", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db2350_0 .net "temp_a_and_out", 0 0, L_0x5c7c33131ba0;  1 drivers
v0x5c7c32db2500_0 .net "temp_a_out", 0 0, L_0x5c7c33131a40;  1 drivers
v0x5c7c32db25a0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33131db0;  1 drivers
v0x5c7c32db2750_0 .net "temp_b_out", 0 0, L_0x5c7c33131c50;  1 drivers
S_0x5c7c32da8570 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32da8390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32da9630_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32da96d0_0 .net "in_b", 0 0, L_0x5c7c33131a40;  alias, 1 drivers
v0x5c7c32da97c0_0 .net "out", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
v0x5c7c32da98e0_0 .net "temp_out", 0 0, L_0x5c7c33131af0;  1 drivers
S_0x5c7c32da87e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32da8570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131af0 .functor NAND 1, L_0x5c7c33133d60, L_0x5c7c33131a40, C4<1>, C4<1>;
v0x5c7c32da8a50_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32da8b60_0 .net "in_b", 0 0, L_0x5c7c33131a40;  alias, 1 drivers
v0x5c7c32da8c20_0 .net "out", 0 0, L_0x5c7c33131af0;  alias, 1 drivers
S_0x5c7c32da8d40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32da8570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32da9480_0 .net "in_a", 0 0, L_0x5c7c33131af0;  alias, 1 drivers
v0x5c7c32da9520_0 .net "out", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
S_0x5c7c32da8f60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32da8d40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131ba0 .functor NAND 1, L_0x5c7c33131af0, L_0x5c7c33131af0, C4<1>, C4<1>;
v0x5c7c32da91d0_0 .net "in_a", 0 0, L_0x5c7c33131af0;  alias, 1 drivers
v0x5c7c32da9290_0 .net "in_b", 0 0, L_0x5c7c33131af0;  alias, 1 drivers
v0x5c7c32da9380_0 .net "out", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
S_0x5c7c32da99a0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32da8390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32daa9d0_0 .net "in_a", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32daaa70_0 .net "in_b", 0 0, L_0x5c7c33131c50;  alias, 1 drivers
v0x5c7c32daab60_0 .net "out", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
v0x5c7c32daac80_0 .net "temp_out", 0 0, L_0x5c7c33131d00;  1 drivers
S_0x5c7c32da9b80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32da99a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131d00 .functor NAND 1, L_0x5c7c33133e00, L_0x5c7c33131c50, C4<1>, C4<1>;
v0x5c7c32da9df0_0 .net "in_a", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32da9f00_0 .net "in_b", 0 0, L_0x5c7c33131c50;  alias, 1 drivers
v0x5c7c32da9fc0_0 .net "out", 0 0, L_0x5c7c33131d00;  alias, 1 drivers
S_0x5c7c32daa0e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32da99a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32daa820_0 .net "in_a", 0 0, L_0x5c7c33131d00;  alias, 1 drivers
v0x5c7c32daa8c0_0 .net "out", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
S_0x5c7c32daa300 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32daa0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131db0 .functor NAND 1, L_0x5c7c33131d00, L_0x5c7c33131d00, C4<1>, C4<1>;
v0x5c7c32daa570_0 .net "in_a", 0 0, L_0x5c7c33131d00;  alias, 1 drivers
v0x5c7c32daa630_0 .net "in_b", 0 0, L_0x5c7c33131d00;  alias, 1 drivers
v0x5c7c32daa720_0 .net "out", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
S_0x5c7c32daadd0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32da8390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dab510_0 .net "in_a", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32dab5b0_0 .net "out", 0 0, L_0x5c7c33131a40;  alias, 1 drivers
S_0x5c7c32daafa0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32daadd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131a40 .functor NAND 1, L_0x5c7c33133e00, L_0x5c7c33133e00, C4<1>, C4<1>;
v0x5c7c32dab1f0_0 .net "in_a", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32dab340_0 .net "in_b", 0 0, L_0x5c7c33133e00;  alias, 1 drivers
v0x5c7c32dab400_0 .net "out", 0 0, L_0x5c7c33131a40;  alias, 1 drivers
S_0x5c7c32dab6b0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32da8390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dabe30_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32dabed0_0 .net "out", 0 0, L_0x5c7c33131c50;  alias, 1 drivers
S_0x5c7c32dab8d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dab6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131c50 .functor NAND 1, L_0x5c7c33133d60, L_0x5c7c33133d60, C4<1>, C4<1>;
v0x5c7c32dabb40_0 .net "in_a", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32dabc90_0 .net "in_b", 0 0, L_0x5c7c33133d60;  alias, 1 drivers
v0x5c7c32dabd50_0 .net "out", 0 0, L_0x5c7c33131c50;  alias, 1 drivers
S_0x5c7c32dabfd0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32da8390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32db1aa0_0 .net "branch1_out", 0 0, L_0x5c7c33131fc0;  1 drivers
v0x5c7c32db1bd0_0 .net "branch2_out", 0 0, L_0x5c7c33132250;  1 drivers
v0x5c7c32db1d20_0 .net "in_a", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
v0x5c7c32db1df0_0 .net "in_b", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
v0x5c7c32db1e90_0 .net "out", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db1f30_0 .net "temp1_out", 0 0, L_0x5c7c33131f10;  1 drivers
v0x5c7c32db1fd0_0 .net "temp2_out", 0 0, L_0x5c7c331321a0;  1 drivers
v0x5c7c32db2070_0 .net "temp3_out", 0 0, L_0x5c7c33132430;  1 drivers
S_0x5c7c32dac250 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32dabfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dad2e0_0 .net "in_a", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
v0x5c7c32dad380_0 .net "in_b", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
v0x5c7c32dad440_0 .net "out", 0 0, L_0x5c7c33131f10;  alias, 1 drivers
v0x5c7c32dad560_0 .net "temp_out", 0 0, L_0x5c7c33131e60;  1 drivers
S_0x5c7c32dac4c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dac250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131e60 .functor NAND 1, L_0x5c7c33131ba0, L_0x5c7c33131ba0, C4<1>, C4<1>;
v0x5c7c32dac730_0 .net "in_a", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
v0x5c7c32dac7f0_0 .net "in_b", 0 0, L_0x5c7c33131ba0;  alias, 1 drivers
v0x5c7c32dac940_0 .net "out", 0 0, L_0x5c7c33131e60;  alias, 1 drivers
S_0x5c7c32daca40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dac250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dad130_0 .net "in_a", 0 0, L_0x5c7c33131e60;  alias, 1 drivers
v0x5c7c32dad1d0_0 .net "out", 0 0, L_0x5c7c33131f10;  alias, 1 drivers
S_0x5c7c32dacc10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32daca40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131f10 .functor NAND 1, L_0x5c7c33131e60, L_0x5c7c33131e60, C4<1>, C4<1>;
v0x5c7c32dace80_0 .net "in_a", 0 0, L_0x5c7c33131e60;  alias, 1 drivers
v0x5c7c32dacf40_0 .net "in_b", 0 0, L_0x5c7c33131e60;  alias, 1 drivers
v0x5c7c32dad030_0 .net "out", 0 0, L_0x5c7c33131f10;  alias, 1 drivers
S_0x5c7c32dad6d0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32dabfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dae700_0 .net "in_a", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
v0x5c7c32dae7a0_0 .net "in_b", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
v0x5c7c32dae860_0 .net "out", 0 0, L_0x5c7c331321a0;  alias, 1 drivers
v0x5c7c32dae980_0 .net "temp_out", 0 0, L_0x5c7c32db0520;  1 drivers
S_0x5c7c32dad8b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dad6d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32db0520 .functor NAND 1, L_0x5c7c33131db0, L_0x5c7c33131db0, C4<1>, C4<1>;
v0x5c7c32dadb20_0 .net "in_a", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
v0x5c7c32dadbe0_0 .net "in_b", 0 0, L_0x5c7c33131db0;  alias, 1 drivers
v0x5c7c32dadd30_0 .net "out", 0 0, L_0x5c7c32db0520;  alias, 1 drivers
S_0x5c7c32dade30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dad6d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dae550_0 .net "in_a", 0 0, L_0x5c7c32db0520;  alias, 1 drivers
v0x5c7c32dae5f0_0 .net "out", 0 0, L_0x5c7c331321a0;  alias, 1 drivers
S_0x5c7c32dae000 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dade30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331321a0 .functor NAND 1, L_0x5c7c32db0520, L_0x5c7c32db0520, C4<1>, C4<1>;
v0x5c7c32dae270_0 .net "in_a", 0 0, L_0x5c7c32db0520;  alias, 1 drivers
v0x5c7c32dae360_0 .net "in_b", 0 0, L_0x5c7c32db0520;  alias, 1 drivers
v0x5c7c32dae450_0 .net "out", 0 0, L_0x5c7c331321a0;  alias, 1 drivers
S_0x5c7c32daeaf0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32dabfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dafb30_0 .net "in_a", 0 0, L_0x5c7c33131fc0;  alias, 1 drivers
v0x5c7c32dafc00_0 .net "in_b", 0 0, L_0x5c7c33132250;  alias, 1 drivers
v0x5c7c32dafcd0_0 .net "out", 0 0, L_0x5c7c33132430;  alias, 1 drivers
v0x5c7c32dafdf0_0 .net "temp_out", 0 0, L_0x5c7c32db0e90;  1 drivers
S_0x5c7c32daecd0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32daeaf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32db0e90 .functor NAND 1, L_0x5c7c33131fc0, L_0x5c7c33132250, C4<1>, C4<1>;
v0x5c7c32daef20_0 .net "in_a", 0 0, L_0x5c7c33131fc0;  alias, 1 drivers
v0x5c7c32daf000_0 .net "in_b", 0 0, L_0x5c7c33132250;  alias, 1 drivers
v0x5c7c32daf0c0_0 .net "out", 0 0, L_0x5c7c32db0e90;  alias, 1 drivers
S_0x5c7c32daf210 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32daeaf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32daf980_0 .net "in_a", 0 0, L_0x5c7c32db0e90;  alias, 1 drivers
v0x5c7c32dafa20_0 .net "out", 0 0, L_0x5c7c33132430;  alias, 1 drivers
S_0x5c7c32daf430 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32daf210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132430 .functor NAND 1, L_0x5c7c32db0e90, L_0x5c7c32db0e90, C4<1>, C4<1>;
v0x5c7c32daf6a0_0 .net "in_a", 0 0, L_0x5c7c32db0e90;  alias, 1 drivers
v0x5c7c32daf790_0 .net "in_b", 0 0, L_0x5c7c32db0e90;  alias, 1 drivers
v0x5c7c32daf880_0 .net "out", 0 0, L_0x5c7c33132430;  alias, 1 drivers
S_0x5c7c32daff40 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32dabfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db0670_0 .net "in_a", 0 0, L_0x5c7c33131f10;  alias, 1 drivers
v0x5c7c32db0710_0 .net "out", 0 0, L_0x5c7c33131fc0;  alias, 1 drivers
S_0x5c7c32db0110 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32daff40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33131fc0 .functor NAND 1, L_0x5c7c33131f10, L_0x5c7c33131f10, C4<1>, C4<1>;
v0x5c7c32db0380_0 .net "in_a", 0 0, L_0x5c7c33131f10;  alias, 1 drivers
v0x5c7c32db0440_0 .net "in_b", 0 0, L_0x5c7c33131f10;  alias, 1 drivers
v0x5c7c32db0590_0 .net "out", 0 0, L_0x5c7c33131fc0;  alias, 1 drivers
S_0x5c7c32db0810 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32dabfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db0fe0_0 .net "in_a", 0 0, L_0x5c7c331321a0;  alias, 1 drivers
v0x5c7c32db1080_0 .net "out", 0 0, L_0x5c7c33132250;  alias, 1 drivers
S_0x5c7c32db0a80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db0810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132250 .functor NAND 1, L_0x5c7c331321a0, L_0x5c7c331321a0, C4<1>, C4<1>;
v0x5c7c32db0cf0_0 .net "in_a", 0 0, L_0x5c7c331321a0;  alias, 1 drivers
v0x5c7c32db0db0_0 .net "in_b", 0 0, L_0x5c7c331321a0;  alias, 1 drivers
v0x5c7c32db0f00_0 .net "out", 0 0, L_0x5c7c33132250;  alias, 1 drivers
S_0x5c7c32db1180 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32dabfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db1920_0 .net "in_a", 0 0, L_0x5c7c33132430;  alias, 1 drivers
v0x5c7c32db19c0_0 .net "out", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
S_0x5c7c32db13a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db1180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331324e0 .functor NAND 1, L_0x5c7c33132430, L_0x5c7c33132430, C4<1>, C4<1>;
v0x5c7c32db1610_0 .net "in_a", 0 0, L_0x5c7c33132430;  alias, 1 drivers
v0x5c7c32db16d0_0 .net "in_b", 0 0, L_0x5c7c33132430;  alias, 1 drivers
v0x5c7c32db1820_0 .net "out", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
S_0x5c7c32db2d30 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32da6ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32dbe850_0 .net "a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32dbe8f0_0 .net "b", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32dbe9b0_0 .net "carry", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32dbea50_0 .net "sum", 0 0, L_0x5c7c33133410;  alias, 1 drivers
S_0x5c7c32db2f50 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32db2d30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32db3ef0_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db3f90_0 .net "in_b", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db4050_0 .net "out", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32db4170_0 .net "temp_out", 0 0, L_0x5c7c32db17b0;  1 drivers
S_0x5c7c32db3100 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32db2f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32db17b0 .functor NAND 1, L_0x5c7c331324e0, L_0x5c7c33131580, C4<1>, C4<1>;
v0x5c7c32db3370_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db3430_0 .net "in_b", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db34f0_0 .net "out", 0 0, L_0x5c7c32db17b0;  alias, 1 drivers
S_0x5c7c32db3620 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32db2f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db3d40_0 .net "in_a", 0 0, L_0x5c7c32db17b0;  alias, 1 drivers
v0x5c7c32db3de0_0 .net "out", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
S_0x5c7c32db37f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db3620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132ae0 .functor NAND 1, L_0x5c7c32db17b0, L_0x5c7c32db17b0, C4<1>, C4<1>;
v0x5c7c32db3a60_0 .net "in_a", 0 0, L_0x5c7c32db17b0;  alias, 1 drivers
v0x5c7c32db3b50_0 .net "in_b", 0 0, L_0x5c7c32db17b0;  alias, 1 drivers
v0x5c7c32db3c40_0 .net "out", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
S_0x5c7c32db42e0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32db2d30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dbe170_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32dbe210_0 .net "in_b", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32dbe2d0_0 .net "out", 0 0, L_0x5c7c33133410;  alias, 1 drivers
v0x5c7c32dbe370_0 .net "temp_a_and_out", 0 0, L_0x5c7c33132cf0;  1 drivers
v0x5c7c32dbe520_0 .net "temp_a_out", 0 0, L_0x5c7c33132b90;  1 drivers
v0x5c7c32dbe5c0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33132f00;  1 drivers
v0x5c7c32dbe770_0 .net "temp_b_out", 0 0, L_0x5c7c33132da0;  1 drivers
S_0x5c7c32db44c0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32db42e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32db5560_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db5710_0 .net "in_b", 0 0, L_0x5c7c33132b90;  alias, 1 drivers
v0x5c7c32db5800_0 .net "out", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
v0x5c7c32db5920_0 .net "temp_out", 0 0, L_0x5c7c33132c40;  1 drivers
S_0x5c7c32db4730 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32db44c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132c40 .functor NAND 1, L_0x5c7c331324e0, L_0x5c7c33132b90, C4<1>, C4<1>;
v0x5c7c32db49a0_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db4a60_0 .net "in_b", 0 0, L_0x5c7c33132b90;  alias, 1 drivers
v0x5c7c32db4b20_0 .net "out", 0 0, L_0x5c7c33132c40;  alias, 1 drivers
S_0x5c7c32db4c40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32db44c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db53b0_0 .net "in_a", 0 0, L_0x5c7c33132c40;  alias, 1 drivers
v0x5c7c32db5450_0 .net "out", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
S_0x5c7c32db4e60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db4c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132cf0 .functor NAND 1, L_0x5c7c33132c40, L_0x5c7c33132c40, C4<1>, C4<1>;
v0x5c7c32db50d0_0 .net "in_a", 0 0, L_0x5c7c33132c40;  alias, 1 drivers
v0x5c7c32db51c0_0 .net "in_b", 0 0, L_0x5c7c33132c40;  alias, 1 drivers
v0x5c7c32db52b0_0 .net "out", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
S_0x5c7c32db59e0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32db42e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32db69f0_0 .net "in_a", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db6a90_0 .net "in_b", 0 0, L_0x5c7c33132da0;  alias, 1 drivers
v0x5c7c32db6b80_0 .net "out", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
v0x5c7c32db6ca0_0 .net "temp_out", 0 0, L_0x5c7c33132e50;  1 drivers
S_0x5c7c32db5bc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32db59e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132e50 .functor NAND 1, L_0x5c7c33131580, L_0x5c7c33132da0, C4<1>, C4<1>;
v0x5c7c32db5e30_0 .net "in_a", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db5ef0_0 .net "in_b", 0 0, L_0x5c7c33132da0;  alias, 1 drivers
v0x5c7c32db5fb0_0 .net "out", 0 0, L_0x5c7c33132e50;  alias, 1 drivers
S_0x5c7c32db60d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32db59e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db6840_0 .net "in_a", 0 0, L_0x5c7c33132e50;  alias, 1 drivers
v0x5c7c32db68e0_0 .net "out", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
S_0x5c7c32db62f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db60d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132f00 .functor NAND 1, L_0x5c7c33132e50, L_0x5c7c33132e50, C4<1>, C4<1>;
v0x5c7c32db6560_0 .net "in_a", 0 0, L_0x5c7c33132e50;  alias, 1 drivers
v0x5c7c32db6650_0 .net "in_b", 0 0, L_0x5c7c33132e50;  alias, 1 drivers
v0x5c7c32db6740_0 .net "out", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
S_0x5c7c32db6df0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32db42e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db7600_0 .net "in_a", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db76a0_0 .net "out", 0 0, L_0x5c7c33132b90;  alias, 1 drivers
S_0x5c7c32db6fc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db6df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132b90 .functor NAND 1, L_0x5c7c33131580, L_0x5c7c33131580, C4<1>, C4<1>;
v0x5c7c32db7210_0 .net "in_a", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db73e0_0 .net "in_b", 0 0, L_0x5c7c33131580;  alias, 1 drivers
v0x5c7c32db74a0_0 .net "out", 0 0, L_0x5c7c33132b90;  alias, 1 drivers
S_0x5c7c32db77a0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32db42e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db7ee0_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db7f80_0 .net "out", 0 0, L_0x5c7c33132da0;  alias, 1 drivers
S_0x5c7c32db79c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db77a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132da0 .functor NAND 1, L_0x5c7c331324e0, L_0x5c7c331324e0, C4<1>, C4<1>;
v0x5c7c32db7c30_0 .net "in_a", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db7cf0_0 .net "in_b", 0 0, L_0x5c7c331324e0;  alias, 1 drivers
v0x5c7c32db7db0_0 .net "out", 0 0, L_0x5c7c33132da0;  alias, 1 drivers
S_0x5c7c32db8080 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32db42e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dbdac0_0 .net "branch1_out", 0 0, L_0x5c7c33133110;  1 drivers
v0x5c7c32dbdbf0_0 .net "branch2_out", 0 0, L_0x5c7c33133290;  1 drivers
v0x5c7c32dbdd40_0 .net "in_a", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
v0x5c7c32dbde10_0 .net "in_b", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
v0x5c7c32dbdeb0_0 .net "out", 0 0, L_0x5c7c33133410;  alias, 1 drivers
v0x5c7c32dbdf50_0 .net "temp1_out", 0 0, L_0x5c7c33133060;  1 drivers
v0x5c7c32dbdff0_0 .net "temp2_out", 0 0, L_0x5c7c331331e0;  1 drivers
v0x5c7c32dbe090_0 .net "temp3_out", 0 0, L_0x5c7c33133360;  1 drivers
S_0x5c7c32db8300 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32db8080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32db9300_0 .net "in_a", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
v0x5c7c32db93a0_0 .net "in_b", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
v0x5c7c32db9460_0 .net "out", 0 0, L_0x5c7c33133060;  alias, 1 drivers
v0x5c7c32db9580_0 .net "temp_out", 0 0, L_0x5c7c33132fb0;  1 drivers
S_0x5c7c32db8570 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32db8300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33132fb0 .functor NAND 1, L_0x5c7c33132cf0, L_0x5c7c33132cf0, C4<1>, C4<1>;
v0x5c7c32db87e0_0 .net "in_a", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
v0x5c7c32db88a0_0 .net "in_b", 0 0, L_0x5c7c33132cf0;  alias, 1 drivers
v0x5c7c32db8960_0 .net "out", 0 0, L_0x5c7c33132fb0;  alias, 1 drivers
S_0x5c7c32db8a60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32db8300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32db9150_0 .net "in_a", 0 0, L_0x5c7c33132fb0;  alias, 1 drivers
v0x5c7c32db91f0_0 .net "out", 0 0, L_0x5c7c33133060;  alias, 1 drivers
S_0x5c7c32db8c30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db8a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133060 .functor NAND 1, L_0x5c7c33132fb0, L_0x5c7c33132fb0, C4<1>, C4<1>;
v0x5c7c32db8ea0_0 .net "in_a", 0 0, L_0x5c7c33132fb0;  alias, 1 drivers
v0x5c7c32db8f60_0 .net "in_b", 0 0, L_0x5c7c33132fb0;  alias, 1 drivers
v0x5c7c32db9050_0 .net "out", 0 0, L_0x5c7c33133060;  alias, 1 drivers
S_0x5c7c32db96f0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32db8080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dba720_0 .net "in_a", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
v0x5c7c32dba7c0_0 .net "in_b", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
v0x5c7c32dba880_0 .net "out", 0 0, L_0x5c7c331331e0;  alias, 1 drivers
v0x5c7c32dba9a0_0 .net "temp_out", 0 0, L_0x5c7c32dbc540;  1 drivers
S_0x5c7c32db98d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32db96f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dbc540 .functor NAND 1, L_0x5c7c33132f00, L_0x5c7c33132f00, C4<1>, C4<1>;
v0x5c7c32db9b40_0 .net "in_a", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
v0x5c7c32db9c00_0 .net "in_b", 0 0, L_0x5c7c33132f00;  alias, 1 drivers
v0x5c7c32db9d50_0 .net "out", 0 0, L_0x5c7c32dbc540;  alias, 1 drivers
S_0x5c7c32db9e50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32db96f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dba570_0 .net "in_a", 0 0, L_0x5c7c32dbc540;  alias, 1 drivers
v0x5c7c32dba610_0 .net "out", 0 0, L_0x5c7c331331e0;  alias, 1 drivers
S_0x5c7c32dba020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32db9e50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331331e0 .functor NAND 1, L_0x5c7c32dbc540, L_0x5c7c32dbc540, C4<1>, C4<1>;
v0x5c7c32dba290_0 .net "in_a", 0 0, L_0x5c7c32dbc540;  alias, 1 drivers
v0x5c7c32dba380_0 .net "in_b", 0 0, L_0x5c7c32dbc540;  alias, 1 drivers
v0x5c7c32dba470_0 .net "out", 0 0, L_0x5c7c331331e0;  alias, 1 drivers
S_0x5c7c32dbab10 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32db8080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dbbb50_0 .net "in_a", 0 0, L_0x5c7c33133110;  alias, 1 drivers
v0x5c7c32dbbc20_0 .net "in_b", 0 0, L_0x5c7c33133290;  alias, 1 drivers
v0x5c7c32dbbcf0_0 .net "out", 0 0, L_0x5c7c33133360;  alias, 1 drivers
v0x5c7c32dbbe10_0 .net "temp_out", 0 0, L_0x5c7c32dbceb0;  1 drivers
S_0x5c7c32dbacf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dbab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dbceb0 .functor NAND 1, L_0x5c7c33133110, L_0x5c7c33133290, C4<1>, C4<1>;
v0x5c7c32dbaf40_0 .net "in_a", 0 0, L_0x5c7c33133110;  alias, 1 drivers
v0x5c7c32dbb020_0 .net "in_b", 0 0, L_0x5c7c33133290;  alias, 1 drivers
v0x5c7c32dbb0e0_0 .net "out", 0 0, L_0x5c7c32dbceb0;  alias, 1 drivers
S_0x5c7c32dbb230 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dbab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dbb9a0_0 .net "in_a", 0 0, L_0x5c7c32dbceb0;  alias, 1 drivers
v0x5c7c32dbba40_0 .net "out", 0 0, L_0x5c7c33133360;  alias, 1 drivers
S_0x5c7c32dbb450 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dbb230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133360 .functor NAND 1, L_0x5c7c32dbceb0, L_0x5c7c32dbceb0, C4<1>, C4<1>;
v0x5c7c32dbb6c0_0 .net "in_a", 0 0, L_0x5c7c32dbceb0;  alias, 1 drivers
v0x5c7c32dbb7b0_0 .net "in_b", 0 0, L_0x5c7c32dbceb0;  alias, 1 drivers
v0x5c7c32dbb8a0_0 .net "out", 0 0, L_0x5c7c33133360;  alias, 1 drivers
S_0x5c7c32dbbf60 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32db8080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dbc690_0 .net "in_a", 0 0, L_0x5c7c33133060;  alias, 1 drivers
v0x5c7c32dbc730_0 .net "out", 0 0, L_0x5c7c33133110;  alias, 1 drivers
S_0x5c7c32dbc130 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dbbf60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133110 .functor NAND 1, L_0x5c7c33133060, L_0x5c7c33133060, C4<1>, C4<1>;
v0x5c7c32dbc3a0_0 .net "in_a", 0 0, L_0x5c7c33133060;  alias, 1 drivers
v0x5c7c32dbc460_0 .net "in_b", 0 0, L_0x5c7c33133060;  alias, 1 drivers
v0x5c7c32dbc5b0_0 .net "out", 0 0, L_0x5c7c33133110;  alias, 1 drivers
S_0x5c7c32dbc830 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32db8080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dbd000_0 .net "in_a", 0 0, L_0x5c7c331331e0;  alias, 1 drivers
v0x5c7c32dbd0a0_0 .net "out", 0 0, L_0x5c7c33133290;  alias, 1 drivers
S_0x5c7c32dbcaa0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dbc830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133290 .functor NAND 1, L_0x5c7c331331e0, L_0x5c7c331331e0, C4<1>, C4<1>;
v0x5c7c32dbcd10_0 .net "in_a", 0 0, L_0x5c7c331331e0;  alias, 1 drivers
v0x5c7c32dbcdd0_0 .net "in_b", 0 0, L_0x5c7c331331e0;  alias, 1 drivers
v0x5c7c32dbcf20_0 .net "out", 0 0, L_0x5c7c33133290;  alias, 1 drivers
S_0x5c7c32dbd1a0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32db8080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dbd940_0 .net "in_a", 0 0, L_0x5c7c33133360;  alias, 1 drivers
v0x5c7c32dbd9e0_0 .net "out", 0 0, L_0x5c7c33133410;  alias, 1 drivers
S_0x5c7c32dbd3c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dbd1a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133410 .functor NAND 1, L_0x5c7c33133360, L_0x5c7c33133360, C4<1>, C4<1>;
v0x5c7c32dbd630_0 .net "in_a", 0 0, L_0x5c7c33133360;  alias, 1 drivers
v0x5c7c32dbd6f0_0 .net "in_b", 0 0, L_0x5c7c33133360;  alias, 1 drivers
v0x5c7c32dbd840_0 .net "out", 0 0, L_0x5c7c33133410;  alias, 1 drivers
S_0x5c7c32dbebc0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32da6ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dc45b0_0 .net "branch1_out", 0 0, L_0x5c7c331336a0;  1 drivers
v0x5c7c32dc46e0_0 .net "branch2_out", 0 0, L_0x5c7c33133930;  1 drivers
v0x5c7c32dc4830_0 .net "in_a", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32dc4a10_0 .net "in_b", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32dc4bc0_0 .net "out", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dc4c60_0 .net "temp1_out", 0 0, L_0x5c7c331335f0;  1 drivers
v0x5c7c32dc4d00_0 .net "temp2_out", 0 0, L_0x5c7c33133880;  1 drivers
v0x5c7c32dc4da0_0 .net "temp3_out", 0 0, L_0x5c7c33133b10;  1 drivers
S_0x5c7c32dbed50 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32dbebc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dbfdf0_0 .net "in_a", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32dbfe90_0 .net "in_b", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32dbff50_0 .net "out", 0 0, L_0x5c7c331335f0;  alias, 1 drivers
v0x5c7c32dc0070_0 .net "temp_out", 0 0, L_0x5c7c32dbd7d0;  1 drivers
S_0x5c7c32dbef70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dbed50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dbd7d0 .functor NAND 1, L_0x5c7c33131990, L_0x5c7c33131990, C4<1>, C4<1>;
v0x5c7c32dbf1e0_0 .net "in_a", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32dbf330_0 .net "in_b", 0 0, L_0x5c7c33131990;  alias, 1 drivers
v0x5c7c32dbf3f0_0 .net "out", 0 0, L_0x5c7c32dbd7d0;  alias, 1 drivers
S_0x5c7c32dbf520 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dbed50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dbfc40_0 .net "in_a", 0 0, L_0x5c7c32dbd7d0;  alias, 1 drivers
v0x5c7c32dbfce0_0 .net "out", 0 0, L_0x5c7c331335f0;  alias, 1 drivers
S_0x5c7c32dbf6f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dbf520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331335f0 .functor NAND 1, L_0x5c7c32dbd7d0, L_0x5c7c32dbd7d0, C4<1>, C4<1>;
v0x5c7c32dbf960_0 .net "in_a", 0 0, L_0x5c7c32dbd7d0;  alias, 1 drivers
v0x5c7c32dbfa50_0 .net "in_b", 0 0, L_0x5c7c32dbd7d0;  alias, 1 drivers
v0x5c7c32dbfb40_0 .net "out", 0 0, L_0x5c7c331335f0;  alias, 1 drivers
S_0x5c7c32dc01e0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32dbebc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dc1210_0 .net "in_a", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32dc12b0_0 .net "in_b", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32dc1370_0 .net "out", 0 0, L_0x5c7c33133880;  alias, 1 drivers
v0x5c7c32dc1490_0 .net "temp_out", 0 0, L_0x5c7c32dc3030;  1 drivers
S_0x5c7c32dc03c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dc01e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dc3030 .functor NAND 1, L_0x5c7c33132ae0, L_0x5c7c33132ae0, C4<1>, C4<1>;
v0x5c7c32dc0630_0 .net "in_a", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32dc0780_0 .net "in_b", 0 0, L_0x5c7c33132ae0;  alias, 1 drivers
v0x5c7c32dc0840_0 .net "out", 0 0, L_0x5c7c32dc3030;  alias, 1 drivers
S_0x5c7c32dc0940 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dc01e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc1060_0 .net "in_a", 0 0, L_0x5c7c32dc3030;  alias, 1 drivers
v0x5c7c32dc1100_0 .net "out", 0 0, L_0x5c7c33133880;  alias, 1 drivers
S_0x5c7c32dc0b10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc0940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133880 .functor NAND 1, L_0x5c7c32dc3030, L_0x5c7c32dc3030, C4<1>, C4<1>;
v0x5c7c32dc0d80_0 .net "in_a", 0 0, L_0x5c7c32dc3030;  alias, 1 drivers
v0x5c7c32dc0e70_0 .net "in_b", 0 0, L_0x5c7c32dc3030;  alias, 1 drivers
v0x5c7c32dc0f60_0 .net "out", 0 0, L_0x5c7c33133880;  alias, 1 drivers
S_0x5c7c32dc1600 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32dbebc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dc2640_0 .net "in_a", 0 0, L_0x5c7c331336a0;  alias, 1 drivers
v0x5c7c32dc2710_0 .net "in_b", 0 0, L_0x5c7c33133930;  alias, 1 drivers
v0x5c7c32dc27e0_0 .net "out", 0 0, L_0x5c7c33133b10;  alias, 1 drivers
v0x5c7c32dc2900_0 .net "temp_out", 0 0, L_0x5c7c32dc39a0;  1 drivers
S_0x5c7c32dc17e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dc1600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dc39a0 .functor NAND 1, L_0x5c7c331336a0, L_0x5c7c33133930, C4<1>, C4<1>;
v0x5c7c32dc1a30_0 .net "in_a", 0 0, L_0x5c7c331336a0;  alias, 1 drivers
v0x5c7c32dc1b10_0 .net "in_b", 0 0, L_0x5c7c33133930;  alias, 1 drivers
v0x5c7c32dc1bd0_0 .net "out", 0 0, L_0x5c7c32dc39a0;  alias, 1 drivers
S_0x5c7c32dc1d20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dc1600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc2490_0 .net "in_a", 0 0, L_0x5c7c32dc39a0;  alias, 1 drivers
v0x5c7c32dc2530_0 .net "out", 0 0, L_0x5c7c33133b10;  alias, 1 drivers
S_0x5c7c32dc1f40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc1d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133b10 .functor NAND 1, L_0x5c7c32dc39a0, L_0x5c7c32dc39a0, C4<1>, C4<1>;
v0x5c7c32dc21b0_0 .net "in_a", 0 0, L_0x5c7c32dc39a0;  alias, 1 drivers
v0x5c7c32dc22a0_0 .net "in_b", 0 0, L_0x5c7c32dc39a0;  alias, 1 drivers
v0x5c7c32dc2390_0 .net "out", 0 0, L_0x5c7c33133b10;  alias, 1 drivers
S_0x5c7c32dc2a50 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32dbebc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc3180_0 .net "in_a", 0 0, L_0x5c7c331335f0;  alias, 1 drivers
v0x5c7c32dc3220_0 .net "out", 0 0, L_0x5c7c331336a0;  alias, 1 drivers
S_0x5c7c32dc2c20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc2a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331336a0 .functor NAND 1, L_0x5c7c331335f0, L_0x5c7c331335f0, C4<1>, C4<1>;
v0x5c7c32dc2e90_0 .net "in_a", 0 0, L_0x5c7c331335f0;  alias, 1 drivers
v0x5c7c32dc2f50_0 .net "in_b", 0 0, L_0x5c7c331335f0;  alias, 1 drivers
v0x5c7c32dc30a0_0 .net "out", 0 0, L_0x5c7c331336a0;  alias, 1 drivers
S_0x5c7c32dc3320 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32dbebc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc3af0_0 .net "in_a", 0 0, L_0x5c7c33133880;  alias, 1 drivers
v0x5c7c32dc3b90_0 .net "out", 0 0, L_0x5c7c33133930;  alias, 1 drivers
S_0x5c7c32dc3590 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc3320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133930 .functor NAND 1, L_0x5c7c33133880, L_0x5c7c33133880, C4<1>, C4<1>;
v0x5c7c32dc3800_0 .net "in_a", 0 0, L_0x5c7c33133880;  alias, 1 drivers
v0x5c7c32dc38c0_0 .net "in_b", 0 0, L_0x5c7c33133880;  alias, 1 drivers
v0x5c7c32dc3a10_0 .net "out", 0 0, L_0x5c7c33133930;  alias, 1 drivers
S_0x5c7c32dc3c90 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32dbebc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc4430_0 .net "in_a", 0 0, L_0x5c7c33133b10;  alias, 1 drivers
v0x5c7c32dc44d0_0 .net "out", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
S_0x5c7c32dc3eb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc3c90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133bc0 .functor NAND 1, L_0x5c7c33133b10, L_0x5c7c33133b10, C4<1>, C4<1>;
v0x5c7c32dc4120_0 .net "in_a", 0 0, L_0x5c7c33133b10;  alias, 1 drivers
v0x5c7c32dc41e0_0 .net "in_b", 0 0, L_0x5c7c33133b10;  alias, 1 drivers
v0x5c7c32dc4330_0 .net "out", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
S_0x5c7c32dc5400 .scope module, "fa_gate16" "FullAdder" 2 21, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32de37b0_0 .net "a", 0 0, L_0x5c7c331363b0;  1 drivers
v0x5c7c32de3850_0 .net "b", 0 0, L_0x5c7c33136660;  1 drivers
v0x5c7c32de3910_0 .net "c", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32de39b0_0 .net "carry", 0 0, L_0x5c7c33136210;  alias, 1 drivers
v0x5c7c32de3a50_0 .net "sum", 0 0, L_0x5c7c33135a60;  1 drivers
v0x5c7c32de3af0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33133fe0;  1 drivers
v0x5c7c32de3b90_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33135130;  1 drivers
v0x5c7c32de3c30_0 .net "tmp_sum_out", 0 0, L_0x5c7c33134b30;  1 drivers
S_0x5c7c32dc55e0 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32dc5400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32dd1160_0 .net "a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dd1310_0 .net "b", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dd14e0_0 .net "carry", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32dd1580_0 .net "sum", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
S_0x5c7c32dc5850 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32dc55e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dc6940_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dc6a10_0 .net "in_b", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc6ae0_0 .net "out", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32dc6c00_0 .net "temp_out", 0 0, L_0x5c7c32dc42c0;  1 drivers
S_0x5c7c32dc5ac0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dc5850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dc42c0 .functor NAND 1, L_0x5c7c331363b0, L_0x5c7c33136660, C4<1>, C4<1>;
v0x5c7c32dc5d30_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dc5e10_0 .net "in_b", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc5ed0_0 .net "out", 0 0, L_0x5c7c32dc42c0;  alias, 1 drivers
S_0x5c7c32dc6020 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dc5850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc6790_0 .net "in_a", 0 0, L_0x5c7c32dc42c0;  alias, 1 drivers
v0x5c7c32dc6830_0 .net "out", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
S_0x5c7c32dc6240 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc6020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33133fe0 .functor NAND 1, L_0x5c7c32dc42c0, L_0x5c7c32dc42c0, C4<1>, C4<1>;
v0x5c7c32dc64b0_0 .net "in_a", 0 0, L_0x5c7c32dc42c0;  alias, 1 drivers
v0x5c7c32dc65a0_0 .net "in_b", 0 0, L_0x5c7c32dc42c0;  alias, 1 drivers
v0x5c7c32dc6690_0 .net "out", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
S_0x5c7c32dc6cc0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32dc55e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd0a80_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dd0b20_0 .net "in_b", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dd0be0_0 .net "out", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd0c80_0 .net "temp_a_and_out", 0 0, L_0x5c7c331341f0;  1 drivers
v0x5c7c32dd0e30_0 .net "temp_a_out", 0 0, L_0x5c7c33134090;  1 drivers
v0x5c7c32dd0ed0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33134400;  1 drivers
v0x5c7c32dd1080_0 .net "temp_b_out", 0 0, L_0x5c7c331342a0;  1 drivers
S_0x5c7c32dc6ea0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32dc6cc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dc7f60_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dc8000_0 .net "in_b", 0 0, L_0x5c7c33134090;  alias, 1 drivers
v0x5c7c32dc80f0_0 .net "out", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
v0x5c7c32dc8210_0 .net "temp_out", 0 0, L_0x5c7c33134140;  1 drivers
S_0x5c7c32dc7110 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dc6ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134140 .functor NAND 1, L_0x5c7c331363b0, L_0x5c7c33134090, C4<1>, C4<1>;
v0x5c7c32dc7380_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dc7490_0 .net "in_b", 0 0, L_0x5c7c33134090;  alias, 1 drivers
v0x5c7c32dc7550_0 .net "out", 0 0, L_0x5c7c33134140;  alias, 1 drivers
S_0x5c7c32dc7670 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dc6ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc7db0_0 .net "in_a", 0 0, L_0x5c7c33134140;  alias, 1 drivers
v0x5c7c32dc7e50_0 .net "out", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
S_0x5c7c32dc7890 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc7670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331341f0 .functor NAND 1, L_0x5c7c33134140, L_0x5c7c33134140, C4<1>, C4<1>;
v0x5c7c32dc7b00_0 .net "in_a", 0 0, L_0x5c7c33134140;  alias, 1 drivers
v0x5c7c32dc7bc0_0 .net "in_b", 0 0, L_0x5c7c33134140;  alias, 1 drivers
v0x5c7c32dc7cb0_0 .net "out", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
S_0x5c7c32dc82d0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32dc6cc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dc9300_0 .net "in_a", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc93a0_0 .net "in_b", 0 0, L_0x5c7c331342a0;  alias, 1 drivers
v0x5c7c32dc9490_0 .net "out", 0 0, L_0x5c7c33134400;  alias, 1 drivers
v0x5c7c32dc95b0_0 .net "temp_out", 0 0, L_0x5c7c33134350;  1 drivers
S_0x5c7c32dc84b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dc82d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134350 .functor NAND 1, L_0x5c7c33136660, L_0x5c7c331342a0, C4<1>, C4<1>;
v0x5c7c32dc8720_0 .net "in_a", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc8830_0 .net "in_b", 0 0, L_0x5c7c331342a0;  alias, 1 drivers
v0x5c7c32dc88f0_0 .net "out", 0 0, L_0x5c7c33134350;  alias, 1 drivers
S_0x5c7c32dc8a10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dc82d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc9150_0 .net "in_a", 0 0, L_0x5c7c33134350;  alias, 1 drivers
v0x5c7c32dc91f0_0 .net "out", 0 0, L_0x5c7c33134400;  alias, 1 drivers
S_0x5c7c32dc8c30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc8a10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134400 .functor NAND 1, L_0x5c7c33134350, L_0x5c7c33134350, C4<1>, C4<1>;
v0x5c7c32dc8ea0_0 .net "in_a", 0 0, L_0x5c7c33134350;  alias, 1 drivers
v0x5c7c32dc8f60_0 .net "in_b", 0 0, L_0x5c7c33134350;  alias, 1 drivers
v0x5c7c32dc9050_0 .net "out", 0 0, L_0x5c7c33134400;  alias, 1 drivers
S_0x5c7c32dc9700 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32dc6cc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dc9e40_0 .net "in_a", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc9ee0_0 .net "out", 0 0, L_0x5c7c33134090;  alias, 1 drivers
S_0x5c7c32dc98d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc9700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134090 .functor NAND 1, L_0x5c7c33136660, L_0x5c7c33136660, C4<1>, C4<1>;
v0x5c7c32dc9b20_0 .net "in_a", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc9c70_0 .net "in_b", 0 0, L_0x5c7c33136660;  alias, 1 drivers
v0x5c7c32dc9d30_0 .net "out", 0 0, L_0x5c7c33134090;  alias, 1 drivers
S_0x5c7c32dc9fe0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32dc6cc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dca760_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dca800_0 .net "out", 0 0, L_0x5c7c331342a0;  alias, 1 drivers
S_0x5c7c32dca200 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dc9fe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331342a0 .functor NAND 1, L_0x5c7c331363b0, L_0x5c7c331363b0, C4<1>, C4<1>;
v0x5c7c32dca470_0 .net "in_a", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dca5c0_0 .net "in_b", 0 0, L_0x5c7c331363b0;  alias, 1 drivers
v0x5c7c32dca680_0 .net "out", 0 0, L_0x5c7c331342a0;  alias, 1 drivers
S_0x5c7c32dca900 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32dc6cc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd03d0_0 .net "branch1_out", 0 0, L_0x5c7c33134610;  1 drivers
v0x5c7c32dd0500_0 .net "branch2_out", 0 0, L_0x5c7c331348a0;  1 drivers
v0x5c7c32dd0650_0 .net "in_a", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
v0x5c7c32dd0720_0 .net "in_b", 0 0, L_0x5c7c33134400;  alias, 1 drivers
v0x5c7c32dd07c0_0 .net "out", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd0860_0 .net "temp1_out", 0 0, L_0x5c7c33134560;  1 drivers
v0x5c7c32dd0900_0 .net "temp2_out", 0 0, L_0x5c7c331347f0;  1 drivers
v0x5c7c32dd09a0_0 .net "temp3_out", 0 0, L_0x5c7c33134a80;  1 drivers
S_0x5c7c32dcab80 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32dca900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dcbc10_0 .net "in_a", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
v0x5c7c32dcbcb0_0 .net "in_b", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
v0x5c7c32dcbd70_0 .net "out", 0 0, L_0x5c7c33134560;  alias, 1 drivers
v0x5c7c32dcbe90_0 .net "temp_out", 0 0, L_0x5c7c331344b0;  1 drivers
S_0x5c7c32dcadf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dcab80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331344b0 .functor NAND 1, L_0x5c7c331341f0, L_0x5c7c331341f0, C4<1>, C4<1>;
v0x5c7c32dcb060_0 .net "in_a", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
v0x5c7c32dcb120_0 .net "in_b", 0 0, L_0x5c7c331341f0;  alias, 1 drivers
v0x5c7c32dcb270_0 .net "out", 0 0, L_0x5c7c331344b0;  alias, 1 drivers
S_0x5c7c32dcb370 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dcab80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dcba60_0 .net "in_a", 0 0, L_0x5c7c331344b0;  alias, 1 drivers
v0x5c7c32dcbb00_0 .net "out", 0 0, L_0x5c7c33134560;  alias, 1 drivers
S_0x5c7c32dcb540 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dcb370;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134560 .functor NAND 1, L_0x5c7c331344b0, L_0x5c7c331344b0, C4<1>, C4<1>;
v0x5c7c32dcb7b0_0 .net "in_a", 0 0, L_0x5c7c331344b0;  alias, 1 drivers
v0x5c7c32dcb870_0 .net "in_b", 0 0, L_0x5c7c331344b0;  alias, 1 drivers
v0x5c7c32dcb960_0 .net "out", 0 0, L_0x5c7c33134560;  alias, 1 drivers
S_0x5c7c32dcc000 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32dca900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dcd030_0 .net "in_a", 0 0, L_0x5c7c33134400;  alias, 1 drivers
v0x5c7c32dcd0d0_0 .net "in_b", 0 0, L_0x5c7c33134400;  alias, 1 drivers
v0x5c7c32dcd190_0 .net "out", 0 0, L_0x5c7c331347f0;  alias, 1 drivers
v0x5c7c32dcd2b0_0 .net "temp_out", 0 0, L_0x5c7c32dcee50;  1 drivers
S_0x5c7c32dcc1e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dcc000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dcee50 .functor NAND 1, L_0x5c7c33134400, L_0x5c7c33134400, C4<1>, C4<1>;
v0x5c7c32dcc450_0 .net "in_a", 0 0, L_0x5c7c33134400;  alias, 1 drivers
v0x5c7c32dcc510_0 .net "in_b", 0 0, L_0x5c7c33134400;  alias, 1 drivers
v0x5c7c32dcc660_0 .net "out", 0 0, L_0x5c7c32dcee50;  alias, 1 drivers
S_0x5c7c32dcc760 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dcc000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dcce80_0 .net "in_a", 0 0, L_0x5c7c32dcee50;  alias, 1 drivers
v0x5c7c32dccf20_0 .net "out", 0 0, L_0x5c7c331347f0;  alias, 1 drivers
S_0x5c7c32dcc930 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dcc760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331347f0 .functor NAND 1, L_0x5c7c32dcee50, L_0x5c7c32dcee50, C4<1>, C4<1>;
v0x5c7c32dccba0_0 .net "in_a", 0 0, L_0x5c7c32dcee50;  alias, 1 drivers
v0x5c7c32dccc90_0 .net "in_b", 0 0, L_0x5c7c32dcee50;  alias, 1 drivers
v0x5c7c32dccd80_0 .net "out", 0 0, L_0x5c7c331347f0;  alias, 1 drivers
S_0x5c7c32dcd420 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32dca900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dce460_0 .net "in_a", 0 0, L_0x5c7c33134610;  alias, 1 drivers
v0x5c7c32dce530_0 .net "in_b", 0 0, L_0x5c7c331348a0;  alias, 1 drivers
v0x5c7c32dce600_0 .net "out", 0 0, L_0x5c7c33134a80;  alias, 1 drivers
v0x5c7c32dce720_0 .net "temp_out", 0 0, L_0x5c7c32dcf7c0;  1 drivers
S_0x5c7c32dcd600 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dcd420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dcf7c0 .functor NAND 1, L_0x5c7c33134610, L_0x5c7c331348a0, C4<1>, C4<1>;
v0x5c7c32dcd850_0 .net "in_a", 0 0, L_0x5c7c33134610;  alias, 1 drivers
v0x5c7c32dcd930_0 .net "in_b", 0 0, L_0x5c7c331348a0;  alias, 1 drivers
v0x5c7c32dcd9f0_0 .net "out", 0 0, L_0x5c7c32dcf7c0;  alias, 1 drivers
S_0x5c7c32dcdb40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dcd420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dce2b0_0 .net "in_a", 0 0, L_0x5c7c32dcf7c0;  alias, 1 drivers
v0x5c7c32dce350_0 .net "out", 0 0, L_0x5c7c33134a80;  alias, 1 drivers
S_0x5c7c32dcdd60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dcdb40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134a80 .functor NAND 1, L_0x5c7c32dcf7c0, L_0x5c7c32dcf7c0, C4<1>, C4<1>;
v0x5c7c32dcdfd0_0 .net "in_a", 0 0, L_0x5c7c32dcf7c0;  alias, 1 drivers
v0x5c7c32dce0c0_0 .net "in_b", 0 0, L_0x5c7c32dcf7c0;  alias, 1 drivers
v0x5c7c32dce1b0_0 .net "out", 0 0, L_0x5c7c33134a80;  alias, 1 drivers
S_0x5c7c32dce870 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32dca900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dcefa0_0 .net "in_a", 0 0, L_0x5c7c33134560;  alias, 1 drivers
v0x5c7c32dcf040_0 .net "out", 0 0, L_0x5c7c33134610;  alias, 1 drivers
S_0x5c7c32dcea40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dce870;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134610 .functor NAND 1, L_0x5c7c33134560, L_0x5c7c33134560, C4<1>, C4<1>;
v0x5c7c32dcecb0_0 .net "in_a", 0 0, L_0x5c7c33134560;  alias, 1 drivers
v0x5c7c32dced70_0 .net "in_b", 0 0, L_0x5c7c33134560;  alias, 1 drivers
v0x5c7c32dceec0_0 .net "out", 0 0, L_0x5c7c33134610;  alias, 1 drivers
S_0x5c7c32dcf140 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32dca900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dcf910_0 .net "in_a", 0 0, L_0x5c7c331347f0;  alias, 1 drivers
v0x5c7c32dcf9b0_0 .net "out", 0 0, L_0x5c7c331348a0;  alias, 1 drivers
S_0x5c7c32dcf3b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dcf140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331348a0 .functor NAND 1, L_0x5c7c331347f0, L_0x5c7c331347f0, C4<1>, C4<1>;
v0x5c7c32dcf620_0 .net "in_a", 0 0, L_0x5c7c331347f0;  alias, 1 drivers
v0x5c7c32dcf6e0_0 .net "in_b", 0 0, L_0x5c7c331347f0;  alias, 1 drivers
v0x5c7c32dcf830_0 .net "out", 0 0, L_0x5c7c331348a0;  alias, 1 drivers
S_0x5c7c32dcfab0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32dca900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd0250_0 .net "in_a", 0 0, L_0x5c7c33134a80;  alias, 1 drivers
v0x5c7c32dd02f0_0 .net "out", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
S_0x5c7c32dcfcd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dcfab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33134b30 .functor NAND 1, L_0x5c7c33134a80, L_0x5c7c33134a80, C4<1>, C4<1>;
v0x5c7c32dcff40_0 .net "in_a", 0 0, L_0x5c7c33134a80;  alias, 1 drivers
v0x5c7c32dd0000_0 .net "in_b", 0 0, L_0x5c7c33134a80;  alias, 1 drivers
v0x5c7c32dd0150_0 .net "out", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
S_0x5c7c32dd1660 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32dc5400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32ddd180_0 .net "a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32ddd220_0 .net "b", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32ddd2e0_0 .net "carry", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32ddd380_0 .net "sum", 0 0, L_0x5c7c33135a60;  alias, 1 drivers
S_0x5c7c32dd1880 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32dd1660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd2820_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd28c0_0 .net "in_b", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd2980_0 .net "out", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32dd2aa0_0 .net "temp_out", 0 0, L_0x5c7c32dd00e0;  1 drivers
S_0x5c7c32dd1a30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dd1880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dd00e0 .functor NAND 1, L_0x5c7c33134b30, L_0x5c7c33133bc0, C4<1>, C4<1>;
v0x5c7c32dd1ca0_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd1d60_0 .net "in_b", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd1e20_0 .net "out", 0 0, L_0x5c7c32dd00e0;  alias, 1 drivers
S_0x5c7c32dd1f50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dd1880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd2670_0 .net "in_a", 0 0, L_0x5c7c32dd00e0;  alias, 1 drivers
v0x5c7c32dd2710_0 .net "out", 0 0, L_0x5c7c33135130;  alias, 1 drivers
S_0x5c7c32dd2120 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd1f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135130 .functor NAND 1, L_0x5c7c32dd00e0, L_0x5c7c32dd00e0, C4<1>, C4<1>;
v0x5c7c32dd2390_0 .net "in_a", 0 0, L_0x5c7c32dd00e0;  alias, 1 drivers
v0x5c7c32dd2480_0 .net "in_b", 0 0, L_0x5c7c32dd00e0;  alias, 1 drivers
v0x5c7c32dd2570_0 .net "out", 0 0, L_0x5c7c33135130;  alias, 1 drivers
S_0x5c7c32dd2c10 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32dd1660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ddcaa0_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32ddcb40_0 .net "in_b", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32ddcc00_0 .net "out", 0 0, L_0x5c7c33135a60;  alias, 1 drivers
v0x5c7c32ddcca0_0 .net "temp_a_and_out", 0 0, L_0x5c7c33135340;  1 drivers
v0x5c7c32ddce50_0 .net "temp_a_out", 0 0, L_0x5c7c331351e0;  1 drivers
v0x5c7c32ddcef0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33135550;  1 drivers
v0x5c7c32ddd0a0_0 .net "temp_b_out", 0 0, L_0x5c7c331353f0;  1 drivers
S_0x5c7c32dd2df0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32dd2c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd3e90_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd4040_0 .net "in_b", 0 0, L_0x5c7c331351e0;  alias, 1 drivers
v0x5c7c32dd4130_0 .net "out", 0 0, L_0x5c7c33135340;  alias, 1 drivers
v0x5c7c32dd4250_0 .net "temp_out", 0 0, L_0x5c7c33135290;  1 drivers
S_0x5c7c32dd3060 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dd2df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135290 .functor NAND 1, L_0x5c7c33134b30, L_0x5c7c331351e0, C4<1>, C4<1>;
v0x5c7c32dd32d0_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd3390_0 .net "in_b", 0 0, L_0x5c7c331351e0;  alias, 1 drivers
v0x5c7c32dd3450_0 .net "out", 0 0, L_0x5c7c33135290;  alias, 1 drivers
S_0x5c7c32dd3570 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dd2df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd3ce0_0 .net "in_a", 0 0, L_0x5c7c33135290;  alias, 1 drivers
v0x5c7c32dd3d80_0 .net "out", 0 0, L_0x5c7c33135340;  alias, 1 drivers
S_0x5c7c32dd3790 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd3570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135340 .functor NAND 1, L_0x5c7c33135290, L_0x5c7c33135290, C4<1>, C4<1>;
v0x5c7c32dd3a00_0 .net "in_a", 0 0, L_0x5c7c33135290;  alias, 1 drivers
v0x5c7c32dd3af0_0 .net "in_b", 0 0, L_0x5c7c33135290;  alias, 1 drivers
v0x5c7c32dd3be0_0 .net "out", 0 0, L_0x5c7c33135340;  alias, 1 drivers
S_0x5c7c32dd4310 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32dd2c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd5320_0 .net "in_a", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd53c0_0 .net "in_b", 0 0, L_0x5c7c331353f0;  alias, 1 drivers
v0x5c7c32dd54b0_0 .net "out", 0 0, L_0x5c7c33135550;  alias, 1 drivers
v0x5c7c32dd55d0_0 .net "temp_out", 0 0, L_0x5c7c331354a0;  1 drivers
S_0x5c7c32dd44f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dd4310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331354a0 .functor NAND 1, L_0x5c7c33133bc0, L_0x5c7c331353f0, C4<1>, C4<1>;
v0x5c7c32dd4760_0 .net "in_a", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd4820_0 .net "in_b", 0 0, L_0x5c7c331353f0;  alias, 1 drivers
v0x5c7c32dd48e0_0 .net "out", 0 0, L_0x5c7c331354a0;  alias, 1 drivers
S_0x5c7c32dd4a00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dd4310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd5170_0 .net "in_a", 0 0, L_0x5c7c331354a0;  alias, 1 drivers
v0x5c7c32dd5210_0 .net "out", 0 0, L_0x5c7c33135550;  alias, 1 drivers
S_0x5c7c32dd4c20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd4a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135550 .functor NAND 1, L_0x5c7c331354a0, L_0x5c7c331354a0, C4<1>, C4<1>;
v0x5c7c32dd4e90_0 .net "in_a", 0 0, L_0x5c7c331354a0;  alias, 1 drivers
v0x5c7c32dd4f80_0 .net "in_b", 0 0, L_0x5c7c331354a0;  alias, 1 drivers
v0x5c7c32dd5070_0 .net "out", 0 0, L_0x5c7c33135550;  alias, 1 drivers
S_0x5c7c32dd5720 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32dd2c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd5f30_0 .net "in_a", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd5fd0_0 .net "out", 0 0, L_0x5c7c331351e0;  alias, 1 drivers
S_0x5c7c32dd58f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd5720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331351e0 .functor NAND 1, L_0x5c7c33133bc0, L_0x5c7c33133bc0, C4<1>, C4<1>;
v0x5c7c32dd5b40_0 .net "in_a", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd5d10_0 .net "in_b", 0 0, L_0x5c7c33133bc0;  alias, 1 drivers
v0x5c7c32dd5dd0_0 .net "out", 0 0, L_0x5c7c331351e0;  alias, 1 drivers
S_0x5c7c32dd60d0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32dd2c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd6810_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd68b0_0 .net "out", 0 0, L_0x5c7c331353f0;  alias, 1 drivers
S_0x5c7c32dd62f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd60d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331353f0 .functor NAND 1, L_0x5c7c33134b30, L_0x5c7c33134b30, C4<1>, C4<1>;
v0x5c7c32dd6560_0 .net "in_a", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd6620_0 .net "in_b", 0 0, L_0x5c7c33134b30;  alias, 1 drivers
v0x5c7c32dd66e0_0 .net "out", 0 0, L_0x5c7c331353f0;  alias, 1 drivers
S_0x5c7c32dd69b0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32dd2c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ddc3f0_0 .net "branch1_out", 0 0, L_0x5c7c33135760;  1 drivers
v0x5c7c32ddc520_0 .net "branch2_out", 0 0, L_0x5c7c331358e0;  1 drivers
v0x5c7c32ddc670_0 .net "in_a", 0 0, L_0x5c7c33135340;  alias, 1 drivers
v0x5c7c32ddc740_0 .net "in_b", 0 0, L_0x5c7c33135550;  alias, 1 drivers
v0x5c7c32ddc7e0_0 .net "out", 0 0, L_0x5c7c33135a60;  alias, 1 drivers
v0x5c7c32ddc880_0 .net "temp1_out", 0 0, L_0x5c7c331356b0;  1 drivers
v0x5c7c32ddc920_0 .net "temp2_out", 0 0, L_0x5c7c33135830;  1 drivers
v0x5c7c32ddc9c0_0 .net "temp3_out", 0 0, L_0x5c7c331359b0;  1 drivers
S_0x5c7c32dd6c30 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32dd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd7c30_0 .net "in_a", 0 0, L_0x5c7c33135340;  alias, 1 drivers
v0x5c7c32dd7cd0_0 .net "in_b", 0 0, L_0x5c7c33135340;  alias, 1 drivers
v0x5c7c32dd7d90_0 .net "out", 0 0, L_0x5c7c331356b0;  alias, 1 drivers
v0x5c7c32dd7eb0_0 .net "temp_out", 0 0, L_0x5c7c33135600;  1 drivers
S_0x5c7c32dd6ea0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dd6c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135600 .functor NAND 1, L_0x5c7c33135340, L_0x5c7c33135340, C4<1>, C4<1>;
v0x5c7c32dd7110_0 .net "in_a", 0 0, L_0x5c7c33135340;  alias, 1 drivers
v0x5c7c32dd71d0_0 .net "in_b", 0 0, L_0x5c7c33135340;  alias, 1 drivers
v0x5c7c32dd7290_0 .net "out", 0 0, L_0x5c7c33135600;  alias, 1 drivers
S_0x5c7c32dd7390 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dd6c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd7a80_0 .net "in_a", 0 0, L_0x5c7c33135600;  alias, 1 drivers
v0x5c7c32dd7b20_0 .net "out", 0 0, L_0x5c7c331356b0;  alias, 1 drivers
S_0x5c7c32dd7560 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd7390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331356b0 .functor NAND 1, L_0x5c7c33135600, L_0x5c7c33135600, C4<1>, C4<1>;
v0x5c7c32dd77d0_0 .net "in_a", 0 0, L_0x5c7c33135600;  alias, 1 drivers
v0x5c7c32dd7890_0 .net "in_b", 0 0, L_0x5c7c33135600;  alias, 1 drivers
v0x5c7c32dd7980_0 .net "out", 0 0, L_0x5c7c331356b0;  alias, 1 drivers
S_0x5c7c32dd8020 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32dd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dd9050_0 .net "in_a", 0 0, L_0x5c7c33135550;  alias, 1 drivers
v0x5c7c32dd90f0_0 .net "in_b", 0 0, L_0x5c7c33135550;  alias, 1 drivers
v0x5c7c32dd91b0_0 .net "out", 0 0, L_0x5c7c33135830;  alias, 1 drivers
v0x5c7c32dd92d0_0 .net "temp_out", 0 0, L_0x5c7c32ddae70;  1 drivers
S_0x5c7c32dd8200 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dd8020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ddae70 .functor NAND 1, L_0x5c7c33135550, L_0x5c7c33135550, C4<1>, C4<1>;
v0x5c7c32dd8470_0 .net "in_a", 0 0, L_0x5c7c33135550;  alias, 1 drivers
v0x5c7c32dd8530_0 .net "in_b", 0 0, L_0x5c7c33135550;  alias, 1 drivers
v0x5c7c32dd8680_0 .net "out", 0 0, L_0x5c7c32ddae70;  alias, 1 drivers
S_0x5c7c32dd8780 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dd8020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dd8ea0_0 .net "in_a", 0 0, L_0x5c7c32ddae70;  alias, 1 drivers
v0x5c7c32dd8f40_0 .net "out", 0 0, L_0x5c7c33135830;  alias, 1 drivers
S_0x5c7c32dd8950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd8780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135830 .functor NAND 1, L_0x5c7c32ddae70, L_0x5c7c32ddae70, C4<1>, C4<1>;
v0x5c7c32dd8bc0_0 .net "in_a", 0 0, L_0x5c7c32ddae70;  alias, 1 drivers
v0x5c7c32dd8cb0_0 .net "in_b", 0 0, L_0x5c7c32ddae70;  alias, 1 drivers
v0x5c7c32dd8da0_0 .net "out", 0 0, L_0x5c7c33135830;  alias, 1 drivers
S_0x5c7c32dd9440 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32dd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dda480_0 .net "in_a", 0 0, L_0x5c7c33135760;  alias, 1 drivers
v0x5c7c32dda550_0 .net "in_b", 0 0, L_0x5c7c331358e0;  alias, 1 drivers
v0x5c7c32dda620_0 .net "out", 0 0, L_0x5c7c331359b0;  alias, 1 drivers
v0x5c7c32dda740_0 .net "temp_out", 0 0, L_0x5c7c32ddb7e0;  1 drivers
S_0x5c7c32dd9620 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dd9440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ddb7e0 .functor NAND 1, L_0x5c7c33135760, L_0x5c7c331358e0, C4<1>, C4<1>;
v0x5c7c32dd9870_0 .net "in_a", 0 0, L_0x5c7c33135760;  alias, 1 drivers
v0x5c7c32dd9950_0 .net "in_b", 0 0, L_0x5c7c331358e0;  alias, 1 drivers
v0x5c7c32dd9a10_0 .net "out", 0 0, L_0x5c7c32ddb7e0;  alias, 1 drivers
S_0x5c7c32dd9b60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dd9440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dda2d0_0 .net "in_a", 0 0, L_0x5c7c32ddb7e0;  alias, 1 drivers
v0x5c7c32dda370_0 .net "out", 0 0, L_0x5c7c331359b0;  alias, 1 drivers
S_0x5c7c32dd9d80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dd9b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331359b0 .functor NAND 1, L_0x5c7c32ddb7e0, L_0x5c7c32ddb7e0, C4<1>, C4<1>;
v0x5c7c32dd9ff0_0 .net "in_a", 0 0, L_0x5c7c32ddb7e0;  alias, 1 drivers
v0x5c7c32dda0e0_0 .net "in_b", 0 0, L_0x5c7c32ddb7e0;  alias, 1 drivers
v0x5c7c32dda1d0_0 .net "out", 0 0, L_0x5c7c331359b0;  alias, 1 drivers
S_0x5c7c32dda890 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32dd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ddafc0_0 .net "in_a", 0 0, L_0x5c7c331356b0;  alias, 1 drivers
v0x5c7c32ddb060_0 .net "out", 0 0, L_0x5c7c33135760;  alias, 1 drivers
S_0x5c7c32ddaa60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dda890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135760 .functor NAND 1, L_0x5c7c331356b0, L_0x5c7c331356b0, C4<1>, C4<1>;
v0x5c7c32ddacd0_0 .net "in_a", 0 0, L_0x5c7c331356b0;  alias, 1 drivers
v0x5c7c32ddad90_0 .net "in_b", 0 0, L_0x5c7c331356b0;  alias, 1 drivers
v0x5c7c32ddaee0_0 .net "out", 0 0, L_0x5c7c33135760;  alias, 1 drivers
S_0x5c7c32ddb160 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32dd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ddb930_0 .net "in_a", 0 0, L_0x5c7c33135830;  alias, 1 drivers
v0x5c7c32ddb9d0_0 .net "out", 0 0, L_0x5c7c331358e0;  alias, 1 drivers
S_0x5c7c32ddb3d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ddb160;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331358e0 .functor NAND 1, L_0x5c7c33135830, L_0x5c7c33135830, C4<1>, C4<1>;
v0x5c7c32ddb640_0 .net "in_a", 0 0, L_0x5c7c33135830;  alias, 1 drivers
v0x5c7c32ddb700_0 .net "in_b", 0 0, L_0x5c7c33135830;  alias, 1 drivers
v0x5c7c32ddb850_0 .net "out", 0 0, L_0x5c7c331358e0;  alias, 1 drivers
S_0x5c7c32ddbad0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32dd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ddc270_0 .net "in_a", 0 0, L_0x5c7c331359b0;  alias, 1 drivers
v0x5c7c32ddc310_0 .net "out", 0 0, L_0x5c7c33135a60;  alias, 1 drivers
S_0x5c7c32ddbcf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ddbad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135a60 .functor NAND 1, L_0x5c7c331359b0, L_0x5c7c331359b0, C4<1>, C4<1>;
v0x5c7c32ddbf60_0 .net "in_a", 0 0, L_0x5c7c331359b0;  alias, 1 drivers
v0x5c7c32ddc020_0 .net "in_b", 0 0, L_0x5c7c331359b0;  alias, 1 drivers
v0x5c7c32ddc170_0 .net "out", 0 0, L_0x5c7c33135a60;  alias, 1 drivers
S_0x5c7c32ddd4f0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32dc5400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32de2ee0_0 .net "branch1_out", 0 0, L_0x5c7c33135cf0;  1 drivers
v0x5c7c32de3010_0 .net "branch2_out", 0 0, L_0x5c7c33135f80;  1 drivers
v0x5c7c32de3160_0 .net "in_a", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32de3340_0 .net "in_b", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32de34f0_0 .net "out", 0 0, L_0x5c7c33136210;  alias, 1 drivers
v0x5c7c32de3590_0 .net "temp1_out", 0 0, L_0x5c7c33135c40;  1 drivers
v0x5c7c32de3630_0 .net "temp2_out", 0 0, L_0x5c7c33135ed0;  1 drivers
v0x5c7c32de36d0_0 .net "temp3_out", 0 0, L_0x5c7c33136160;  1 drivers
S_0x5c7c32ddd680 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32ddd4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dde720_0 .net "in_a", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32dde7c0_0 .net "in_b", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32dde880_0 .net "out", 0 0, L_0x5c7c33135c40;  alias, 1 drivers
v0x5c7c32dde9a0_0 .net "temp_out", 0 0, L_0x5c7c32ddc100;  1 drivers
S_0x5c7c32ddd8a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ddd680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ddc100 .functor NAND 1, L_0x5c7c33133fe0, L_0x5c7c33133fe0, C4<1>, C4<1>;
v0x5c7c32dddb10_0 .net "in_a", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32dddc60_0 .net "in_b", 0 0, L_0x5c7c33133fe0;  alias, 1 drivers
v0x5c7c32dddd20_0 .net "out", 0 0, L_0x5c7c32ddc100;  alias, 1 drivers
S_0x5c7c32ddde50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ddd680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dde570_0 .net "in_a", 0 0, L_0x5c7c32ddc100;  alias, 1 drivers
v0x5c7c32dde610_0 .net "out", 0 0, L_0x5c7c33135c40;  alias, 1 drivers
S_0x5c7c32dde020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ddde50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135c40 .functor NAND 1, L_0x5c7c32ddc100, L_0x5c7c32ddc100, C4<1>, C4<1>;
v0x5c7c32dde290_0 .net "in_a", 0 0, L_0x5c7c32ddc100;  alias, 1 drivers
v0x5c7c32dde380_0 .net "in_b", 0 0, L_0x5c7c32ddc100;  alias, 1 drivers
v0x5c7c32dde470_0 .net "out", 0 0, L_0x5c7c33135c40;  alias, 1 drivers
S_0x5c7c32ddeb10 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32ddd4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ddfb40_0 .net "in_a", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32ddfbe0_0 .net "in_b", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32ddfca0_0 .net "out", 0 0, L_0x5c7c33135ed0;  alias, 1 drivers
v0x5c7c32ddfdc0_0 .net "temp_out", 0 0, L_0x5c7c32de1960;  1 drivers
S_0x5c7c32ddecf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ddeb10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32de1960 .functor NAND 1, L_0x5c7c33135130, L_0x5c7c33135130, C4<1>, C4<1>;
v0x5c7c32ddef60_0 .net "in_a", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32ddf0b0_0 .net "in_b", 0 0, L_0x5c7c33135130;  alias, 1 drivers
v0x5c7c32ddf170_0 .net "out", 0 0, L_0x5c7c32de1960;  alias, 1 drivers
S_0x5c7c32ddf270 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ddeb10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ddf990_0 .net "in_a", 0 0, L_0x5c7c32de1960;  alias, 1 drivers
v0x5c7c32ddfa30_0 .net "out", 0 0, L_0x5c7c33135ed0;  alias, 1 drivers
S_0x5c7c32ddf440 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ddf270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135ed0 .functor NAND 1, L_0x5c7c32de1960, L_0x5c7c32de1960, C4<1>, C4<1>;
v0x5c7c32ddf6b0_0 .net "in_a", 0 0, L_0x5c7c32de1960;  alias, 1 drivers
v0x5c7c32ddf7a0_0 .net "in_b", 0 0, L_0x5c7c32de1960;  alias, 1 drivers
v0x5c7c32ddf890_0 .net "out", 0 0, L_0x5c7c33135ed0;  alias, 1 drivers
S_0x5c7c32ddff30 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32ddd4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32de0f70_0 .net "in_a", 0 0, L_0x5c7c33135cf0;  alias, 1 drivers
v0x5c7c32de1040_0 .net "in_b", 0 0, L_0x5c7c33135f80;  alias, 1 drivers
v0x5c7c32de1110_0 .net "out", 0 0, L_0x5c7c33136160;  alias, 1 drivers
v0x5c7c32de1230_0 .net "temp_out", 0 0, L_0x5c7c32de22d0;  1 drivers
S_0x5c7c32de0110 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ddff30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32de22d0 .functor NAND 1, L_0x5c7c33135cf0, L_0x5c7c33135f80, C4<1>, C4<1>;
v0x5c7c32de0360_0 .net "in_a", 0 0, L_0x5c7c33135cf0;  alias, 1 drivers
v0x5c7c32de0440_0 .net "in_b", 0 0, L_0x5c7c33135f80;  alias, 1 drivers
v0x5c7c32de0500_0 .net "out", 0 0, L_0x5c7c32de22d0;  alias, 1 drivers
S_0x5c7c32de0650 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ddff30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de0dc0_0 .net "in_a", 0 0, L_0x5c7c32de22d0;  alias, 1 drivers
v0x5c7c32de0e60_0 .net "out", 0 0, L_0x5c7c33136160;  alias, 1 drivers
S_0x5c7c32de0870 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de0650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33136160 .functor NAND 1, L_0x5c7c32de22d0, L_0x5c7c32de22d0, C4<1>, C4<1>;
v0x5c7c32de0ae0_0 .net "in_a", 0 0, L_0x5c7c32de22d0;  alias, 1 drivers
v0x5c7c32de0bd0_0 .net "in_b", 0 0, L_0x5c7c32de22d0;  alias, 1 drivers
v0x5c7c32de0cc0_0 .net "out", 0 0, L_0x5c7c33136160;  alias, 1 drivers
S_0x5c7c32de1380 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32ddd4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de1ab0_0 .net "in_a", 0 0, L_0x5c7c33135c40;  alias, 1 drivers
v0x5c7c32de1b50_0 .net "out", 0 0, L_0x5c7c33135cf0;  alias, 1 drivers
S_0x5c7c32de1550 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de1380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135cf0 .functor NAND 1, L_0x5c7c33135c40, L_0x5c7c33135c40, C4<1>, C4<1>;
v0x5c7c32de17c0_0 .net "in_a", 0 0, L_0x5c7c33135c40;  alias, 1 drivers
v0x5c7c32de1880_0 .net "in_b", 0 0, L_0x5c7c33135c40;  alias, 1 drivers
v0x5c7c32de19d0_0 .net "out", 0 0, L_0x5c7c33135cf0;  alias, 1 drivers
S_0x5c7c32de1c50 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32ddd4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de2420_0 .net "in_a", 0 0, L_0x5c7c33135ed0;  alias, 1 drivers
v0x5c7c32de24c0_0 .net "out", 0 0, L_0x5c7c33135f80;  alias, 1 drivers
S_0x5c7c32de1ec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de1c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33135f80 .functor NAND 1, L_0x5c7c33135ed0, L_0x5c7c33135ed0, C4<1>, C4<1>;
v0x5c7c32de2130_0 .net "in_a", 0 0, L_0x5c7c33135ed0;  alias, 1 drivers
v0x5c7c32de21f0_0 .net "in_b", 0 0, L_0x5c7c33135ed0;  alias, 1 drivers
v0x5c7c32de2340_0 .net "out", 0 0, L_0x5c7c33135f80;  alias, 1 drivers
S_0x5c7c32de25c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32ddd4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de2d60_0 .net "in_a", 0 0, L_0x5c7c33136160;  alias, 1 drivers
v0x5c7c32de2e00_0 .net "out", 0 0, L_0x5c7c33136210;  alias, 1 drivers
S_0x5c7c32de27e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de25c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33136210 .functor NAND 1, L_0x5c7c33136160, L_0x5c7c33136160, C4<1>, C4<1>;
v0x5c7c32de2a50_0 .net "in_a", 0 0, L_0x5c7c33136160;  alias, 1 drivers
v0x5c7c32de2b10_0 .net "in_b", 0 0, L_0x5c7c33136160;  alias, 1 drivers
v0x5c7c32de2c60_0 .net "out", 0 0, L_0x5c7c33136210;  alias, 1 drivers
S_0x5c7c32de3d30 .scope module, "fa_gate2" "FullAdder" 2 7, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32e021b0_0 .net "a", 0 0, L_0x5c7c33115020;  1 drivers
v0x5c7c32e02250_0 .net "b", 0 0, L_0x5c7c331150c0;  1 drivers
v0x5c7c32e02310_0 .net "c", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32e023b0_0 .net "carry", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e02450_0 .net "sum", 0 0, L_0x5c7c331146d0;  1 drivers
v0x5c7c32e024f0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33112d40;  1 drivers
v0x5c7c32e02590_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33113da0;  1 drivers
v0x5c7c32e02630_0 .net "tmp_sum_out", 0 0, L_0x5c7c331139b0;  1 drivers
S_0x5c7c32de3f90 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32de3d30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32defb10_0 .net "a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32defcc0_0 .net "b", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32defe90_0 .net "carry", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32deff30_0 .net "sum", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
S_0x5c7c32de4200 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32de3f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32de52f0_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de53c0_0 .net "in_b", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de5490_0 .net "out", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32de55b0_0 .net "temp_out", 0 0, L_0x5c7c33112cb0;  1 drivers
S_0x5c7c32de4470 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32de4200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112cb0 .functor NAND 1, L_0x5c7c33115020, L_0x5c7c331150c0, C4<1>, C4<1>;
v0x5c7c32de46e0_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de47c0_0 .net "in_b", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de4880_0 .net "out", 0 0, L_0x5c7c33112cb0;  alias, 1 drivers
S_0x5c7c32de49d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32de4200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de5140_0 .net "in_a", 0 0, L_0x5c7c33112cb0;  alias, 1 drivers
v0x5c7c32de51e0_0 .net "out", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
S_0x5c7c32de4bf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de49d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112d40 .functor NAND 1, L_0x5c7c33112cb0, L_0x5c7c33112cb0, C4<1>, C4<1>;
v0x5c7c32de4e60_0 .net "in_a", 0 0, L_0x5c7c33112cb0;  alias, 1 drivers
v0x5c7c32de4f50_0 .net "in_b", 0 0, L_0x5c7c33112cb0;  alias, 1 drivers
v0x5c7c32de5040_0 .net "out", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
S_0x5c7c32de5670 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32de3f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32def430_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32def4d0_0 .net "in_b", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32def590_0 .net "out", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32def630_0 .net "temp_a_and_out", 0 0, L_0x5c7c33112f50;  1 drivers
v0x5c7c32def7e0_0 .net "temp_a_out", 0 0, L_0x5c7c33112df0;  1 drivers
v0x5c7c32def880_0 .net "temp_b_and_out", 0 0, L_0x5c7c33113160;  1 drivers
v0x5c7c32defa30_0 .net "temp_b_out", 0 0, L_0x5c7c33113000;  1 drivers
S_0x5c7c32de5850 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32de5670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32de6910_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de69b0_0 .net "in_b", 0 0, L_0x5c7c33112df0;  alias, 1 drivers
v0x5c7c32de6aa0_0 .net "out", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
v0x5c7c32de6bc0_0 .net "temp_out", 0 0, L_0x5c7c33112ea0;  1 drivers
S_0x5c7c32de5ac0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32de5850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112ea0 .functor NAND 1, L_0x5c7c33115020, L_0x5c7c33112df0, C4<1>, C4<1>;
v0x5c7c32de5d30_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de5e40_0 .net "in_b", 0 0, L_0x5c7c33112df0;  alias, 1 drivers
v0x5c7c32de5f00_0 .net "out", 0 0, L_0x5c7c33112ea0;  alias, 1 drivers
S_0x5c7c32de6020 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32de5850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de6760_0 .net "in_a", 0 0, L_0x5c7c33112ea0;  alias, 1 drivers
v0x5c7c32de6800_0 .net "out", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
S_0x5c7c32de6240 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de6020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112f50 .functor NAND 1, L_0x5c7c33112ea0, L_0x5c7c33112ea0, C4<1>, C4<1>;
v0x5c7c32de64b0_0 .net "in_a", 0 0, L_0x5c7c33112ea0;  alias, 1 drivers
v0x5c7c32de6570_0 .net "in_b", 0 0, L_0x5c7c33112ea0;  alias, 1 drivers
v0x5c7c32de6660_0 .net "out", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
S_0x5c7c32de6c80 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32de5670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32de7cb0_0 .net "in_a", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de7d50_0 .net "in_b", 0 0, L_0x5c7c33113000;  alias, 1 drivers
v0x5c7c32de7e40_0 .net "out", 0 0, L_0x5c7c33113160;  alias, 1 drivers
v0x5c7c32de7f60_0 .net "temp_out", 0 0, L_0x5c7c331130b0;  1 drivers
S_0x5c7c32de6e60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32de6c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331130b0 .functor NAND 1, L_0x5c7c331150c0, L_0x5c7c33113000, C4<1>, C4<1>;
v0x5c7c32de70d0_0 .net "in_a", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de71e0_0 .net "in_b", 0 0, L_0x5c7c33113000;  alias, 1 drivers
v0x5c7c32de72a0_0 .net "out", 0 0, L_0x5c7c331130b0;  alias, 1 drivers
S_0x5c7c32de73c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32de6c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de7b00_0 .net "in_a", 0 0, L_0x5c7c331130b0;  alias, 1 drivers
v0x5c7c32de7ba0_0 .net "out", 0 0, L_0x5c7c33113160;  alias, 1 drivers
S_0x5c7c32de75e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de73c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113160 .functor NAND 1, L_0x5c7c331130b0, L_0x5c7c331130b0, C4<1>, C4<1>;
v0x5c7c32de7850_0 .net "in_a", 0 0, L_0x5c7c331130b0;  alias, 1 drivers
v0x5c7c32de7910_0 .net "in_b", 0 0, L_0x5c7c331130b0;  alias, 1 drivers
v0x5c7c32de7a00_0 .net "out", 0 0, L_0x5c7c33113160;  alias, 1 drivers
S_0x5c7c32de80b0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32de5670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de87f0_0 .net "in_a", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de8890_0 .net "out", 0 0, L_0x5c7c33112df0;  alias, 1 drivers
S_0x5c7c32de8280 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de80b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112df0 .functor NAND 1, L_0x5c7c331150c0, L_0x5c7c331150c0, C4<1>, C4<1>;
v0x5c7c32de84d0_0 .net "in_a", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de8620_0 .net "in_b", 0 0, L_0x5c7c331150c0;  alias, 1 drivers
v0x5c7c32de86e0_0 .net "out", 0 0, L_0x5c7c33112df0;  alias, 1 drivers
S_0x5c7c32de8990 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32de5670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32de9110_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de91b0_0 .net "out", 0 0, L_0x5c7c33113000;  alias, 1 drivers
S_0x5c7c32de8bb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de8990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113000 .functor NAND 1, L_0x5c7c33115020, L_0x5c7c33115020, C4<1>, C4<1>;
v0x5c7c32de8e20_0 .net "in_a", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de8f70_0 .net "in_b", 0 0, L_0x5c7c33115020;  alias, 1 drivers
v0x5c7c32de9030_0 .net "out", 0 0, L_0x5c7c33113000;  alias, 1 drivers
S_0x5c7c32de92b0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32de5670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32deed80_0 .net "branch1_out", 0 0, L_0x5c7c33113370;  1 drivers
v0x5c7c32deeeb0_0 .net "branch2_out", 0 0, L_0x5c7c33113690;  1 drivers
v0x5c7c32def000_0 .net "in_a", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
v0x5c7c32def0d0_0 .net "in_b", 0 0, L_0x5c7c33113160;  alias, 1 drivers
v0x5c7c32def170_0 .net "out", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32def210_0 .net "temp1_out", 0 0, L_0x5c7c331132c0;  1 drivers
v0x5c7c32def2b0_0 .net "temp2_out", 0 0, L_0x5c7c331135e0;  1 drivers
v0x5c7c32def350_0 .net "temp3_out", 0 0, L_0x5c7c33113900;  1 drivers
S_0x5c7c32de9530 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32de92b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dea5c0_0 .net "in_a", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
v0x5c7c32dea660_0 .net "in_b", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
v0x5c7c32dea720_0 .net "out", 0 0, L_0x5c7c331132c0;  alias, 1 drivers
v0x5c7c32dea840_0 .net "temp_out", 0 0, L_0x5c7c33113210;  1 drivers
S_0x5c7c32de97a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32de9530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113210 .functor NAND 1, L_0x5c7c33112f50, L_0x5c7c33112f50, C4<1>, C4<1>;
v0x5c7c32de9a10_0 .net "in_a", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
v0x5c7c32de9ad0_0 .net "in_b", 0 0, L_0x5c7c33112f50;  alias, 1 drivers
v0x5c7c32de9c20_0 .net "out", 0 0, L_0x5c7c33113210;  alias, 1 drivers
S_0x5c7c32de9d20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32de9530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dea410_0 .net "in_a", 0 0, L_0x5c7c33113210;  alias, 1 drivers
v0x5c7c32dea4b0_0 .net "out", 0 0, L_0x5c7c331132c0;  alias, 1 drivers
S_0x5c7c32de9ef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32de9d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331132c0 .functor NAND 1, L_0x5c7c33113210, L_0x5c7c33113210, C4<1>, C4<1>;
v0x5c7c32dea160_0 .net "in_a", 0 0, L_0x5c7c33113210;  alias, 1 drivers
v0x5c7c32dea220_0 .net "in_b", 0 0, L_0x5c7c33113210;  alias, 1 drivers
v0x5c7c32dea310_0 .net "out", 0 0, L_0x5c7c331132c0;  alias, 1 drivers
S_0x5c7c32dea9b0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32de92b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32deb9e0_0 .net "in_a", 0 0, L_0x5c7c33113160;  alias, 1 drivers
v0x5c7c32deba80_0 .net "in_b", 0 0, L_0x5c7c33113160;  alias, 1 drivers
v0x5c7c32debb40_0 .net "out", 0 0, L_0x5c7c331135e0;  alias, 1 drivers
v0x5c7c32debc60_0 .net "temp_out", 0 0, L_0x5c7c33113530;  1 drivers
S_0x5c7c32deab90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dea9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113530 .functor NAND 1, L_0x5c7c33113160, L_0x5c7c33113160, C4<1>, C4<1>;
v0x5c7c32deae00_0 .net "in_a", 0 0, L_0x5c7c33113160;  alias, 1 drivers
v0x5c7c32deaec0_0 .net "in_b", 0 0, L_0x5c7c33113160;  alias, 1 drivers
v0x5c7c32deb010_0 .net "out", 0 0, L_0x5c7c33113530;  alias, 1 drivers
S_0x5c7c32deb110 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dea9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32deb830_0 .net "in_a", 0 0, L_0x5c7c33113530;  alias, 1 drivers
v0x5c7c32deb8d0_0 .net "out", 0 0, L_0x5c7c331135e0;  alias, 1 drivers
S_0x5c7c32deb2e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32deb110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331135e0 .functor NAND 1, L_0x5c7c33113530, L_0x5c7c33113530, C4<1>, C4<1>;
v0x5c7c32deb550_0 .net "in_a", 0 0, L_0x5c7c33113530;  alias, 1 drivers
v0x5c7c32deb640_0 .net "in_b", 0 0, L_0x5c7c33113530;  alias, 1 drivers
v0x5c7c32deb730_0 .net "out", 0 0, L_0x5c7c331135e0;  alias, 1 drivers
S_0x5c7c32debdd0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32de92b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dece10_0 .net "in_a", 0 0, L_0x5c7c33113370;  alias, 1 drivers
v0x5c7c32decee0_0 .net "in_b", 0 0, L_0x5c7c33113690;  alias, 1 drivers
v0x5c7c32decfb0_0 .net "out", 0 0, L_0x5c7c33113900;  alias, 1 drivers
v0x5c7c32ded0d0_0 .net "temp_out", 0 0, L_0x5c7c33113850;  1 drivers
S_0x5c7c32debfb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32debdd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113850 .functor NAND 1, L_0x5c7c33113370, L_0x5c7c33113690, C4<1>, C4<1>;
v0x5c7c32dec200_0 .net "in_a", 0 0, L_0x5c7c33113370;  alias, 1 drivers
v0x5c7c32dec2e0_0 .net "in_b", 0 0, L_0x5c7c33113690;  alias, 1 drivers
v0x5c7c32dec3a0_0 .net "out", 0 0, L_0x5c7c33113850;  alias, 1 drivers
S_0x5c7c32dec4f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32debdd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32decc60_0 .net "in_a", 0 0, L_0x5c7c33113850;  alias, 1 drivers
v0x5c7c32decd00_0 .net "out", 0 0, L_0x5c7c33113900;  alias, 1 drivers
S_0x5c7c32dec710 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dec4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113900 .functor NAND 1, L_0x5c7c33113850, L_0x5c7c33113850, C4<1>, C4<1>;
v0x5c7c32dec980_0 .net "in_a", 0 0, L_0x5c7c33113850;  alias, 1 drivers
v0x5c7c32deca70_0 .net "in_b", 0 0, L_0x5c7c33113850;  alias, 1 drivers
v0x5c7c32decb60_0 .net "out", 0 0, L_0x5c7c33113900;  alias, 1 drivers
S_0x5c7c32ded220 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32de92b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ded950_0 .net "in_a", 0 0, L_0x5c7c331132c0;  alias, 1 drivers
v0x5c7c32ded9f0_0 .net "out", 0 0, L_0x5c7c33113370;  alias, 1 drivers
S_0x5c7c32ded3f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ded220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113370 .functor NAND 1, L_0x5c7c331132c0, L_0x5c7c331132c0, C4<1>, C4<1>;
v0x5c7c32ded660_0 .net "in_a", 0 0, L_0x5c7c331132c0;  alias, 1 drivers
v0x5c7c32ded720_0 .net "in_b", 0 0, L_0x5c7c331132c0;  alias, 1 drivers
v0x5c7c32ded870_0 .net "out", 0 0, L_0x5c7c33113370;  alias, 1 drivers
S_0x5c7c32dedaf0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32de92b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dee2c0_0 .net "in_a", 0 0, L_0x5c7c331135e0;  alias, 1 drivers
v0x5c7c32dee360_0 .net "out", 0 0, L_0x5c7c33113690;  alias, 1 drivers
S_0x5c7c32dedd60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dedaf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113690 .functor NAND 1, L_0x5c7c331135e0, L_0x5c7c331135e0, C4<1>, C4<1>;
v0x5c7c32dedfd0_0 .net "in_a", 0 0, L_0x5c7c331135e0;  alias, 1 drivers
v0x5c7c32dee090_0 .net "in_b", 0 0, L_0x5c7c331135e0;  alias, 1 drivers
v0x5c7c32dee1e0_0 .net "out", 0 0, L_0x5c7c33113690;  alias, 1 drivers
S_0x5c7c32dee460 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32de92b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32deec00_0 .net "in_a", 0 0, L_0x5c7c33113900;  alias, 1 drivers
v0x5c7c32deeca0_0 .net "out", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
S_0x5c7c32dee680 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dee460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331139b0 .functor NAND 1, L_0x5c7c33113900, L_0x5c7c33113900, C4<1>, C4<1>;
v0x5c7c32dee8f0_0 .net "in_a", 0 0, L_0x5c7c33113900;  alias, 1 drivers
v0x5c7c32dee9b0_0 .net "in_b", 0 0, L_0x5c7c33113900;  alias, 1 drivers
v0x5c7c32deeb00_0 .net "out", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
S_0x5c7c32df0010 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32de3d30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32dfbb00_0 .net "a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32dfbba0_0 .net "b", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32dfbd70_0 .net "carry", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32dfbe10_0 .net "sum", 0 0, L_0x5c7c331146d0;  alias, 1 drivers
S_0x5c7c32df0230 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32df0010;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32df1240_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df12e0_0 .net "in_b", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df13d0_0 .net "out", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32df14f0_0 .net "temp_out", 0 0, L_0x5c7c32deea90;  1 drivers
S_0x5c7c32df03e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32df0230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32deea90 .functor NAND 1, L_0x5c7c331139b0, L_0x5c7c33111ce0, C4<1>, C4<1>;
v0x5c7c32df0650_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df0710_0 .net "in_b", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df07d0_0 .net "out", 0 0, L_0x5c7c32deea90;  alias, 1 drivers
S_0x5c7c32df0920 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32df0230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df1090_0 .net "in_a", 0 0, L_0x5c7c32deea90;  alias, 1 drivers
v0x5c7c32df1130_0 .net "out", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
S_0x5c7c32df0b40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df0920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113da0 .functor NAND 1, L_0x5c7c32deea90, L_0x5c7c32deea90, C4<1>, C4<1>;
v0x5c7c32df0db0_0 .net "in_a", 0 0, L_0x5c7c32deea90;  alias, 1 drivers
v0x5c7c32df0ea0_0 .net "in_b", 0 0, L_0x5c7c32deea90;  alias, 1 drivers
v0x5c7c32df0f90_0 .net "out", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
S_0x5c7c32df15b0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32df0010;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dfb420_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32dfb4c0_0 .net "in_b", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32dfb580_0 .net "out", 0 0, L_0x5c7c331146d0;  alias, 1 drivers
v0x5c7c32dfb620_0 .net "temp_a_and_out", 0 0, L_0x5c7c33113fb0;  1 drivers
v0x5c7c32dfb7d0_0 .net "temp_a_out", 0 0, L_0x5c7c33113e50;  1 drivers
v0x5c7c32dfb870_0 .net "temp_b_and_out", 0 0, L_0x5c7c331141c0;  1 drivers
v0x5c7c32dfba20_0 .net "temp_b_out", 0 0, L_0x5c7c33114060;  1 drivers
S_0x5c7c32df1790 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32df15b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32df2830_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df29e0_0 .net "in_b", 0 0, L_0x5c7c33113e50;  alias, 1 drivers
v0x5c7c32df2ad0_0 .net "out", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
v0x5c7c32df2bf0_0 .net "temp_out", 0 0, L_0x5c7c33113f00;  1 drivers
S_0x5c7c32df1a00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32df1790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113f00 .functor NAND 1, L_0x5c7c331139b0, L_0x5c7c33113e50, C4<1>, C4<1>;
v0x5c7c32df1c70_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df1d30_0 .net "in_b", 0 0, L_0x5c7c33113e50;  alias, 1 drivers
v0x5c7c32df1df0_0 .net "out", 0 0, L_0x5c7c33113f00;  alias, 1 drivers
S_0x5c7c32df1f10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32df1790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df2680_0 .net "in_a", 0 0, L_0x5c7c33113f00;  alias, 1 drivers
v0x5c7c32df2720_0 .net "out", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
S_0x5c7c32df2130 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df1f10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113fb0 .functor NAND 1, L_0x5c7c33113f00, L_0x5c7c33113f00, C4<1>, C4<1>;
v0x5c7c32df23a0_0 .net "in_a", 0 0, L_0x5c7c33113f00;  alias, 1 drivers
v0x5c7c32df2490_0 .net "in_b", 0 0, L_0x5c7c33113f00;  alias, 1 drivers
v0x5c7c32df2580_0 .net "out", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
S_0x5c7c32df2cb0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32df15b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32df3ce0_0 .net "in_a", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df3d80_0 .net "in_b", 0 0, L_0x5c7c33114060;  alias, 1 drivers
v0x5c7c32df3e70_0 .net "out", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
v0x5c7c32df3f90_0 .net "temp_out", 0 0, L_0x5c7c33114110;  1 drivers
S_0x5c7c32df2e90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32df2cb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114110 .functor NAND 1, L_0x5c7c33111ce0, L_0x5c7c33114060, C4<1>, C4<1>;
v0x5c7c32df3100_0 .net "in_a", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df3210_0 .net "in_b", 0 0, L_0x5c7c33114060;  alias, 1 drivers
v0x5c7c32df32d0_0 .net "out", 0 0, L_0x5c7c33114110;  alias, 1 drivers
S_0x5c7c32df33f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32df2cb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df3b30_0 .net "in_a", 0 0, L_0x5c7c33114110;  alias, 1 drivers
v0x5c7c32df3bd0_0 .net "out", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
S_0x5c7c32df3610 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df33f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331141c0 .functor NAND 1, L_0x5c7c33114110, L_0x5c7c33114110, C4<1>, C4<1>;
v0x5c7c32df3880_0 .net "in_a", 0 0, L_0x5c7c33114110;  alias, 1 drivers
v0x5c7c32df3940_0 .net "in_b", 0 0, L_0x5c7c33114110;  alias, 1 drivers
v0x5c7c32df3a30_0 .net "out", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
S_0x5c7c32df40e0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32df15b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df4820_0 .net "in_a", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df48c0_0 .net "out", 0 0, L_0x5c7c33113e50;  alias, 1 drivers
S_0x5c7c32df42b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df40e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33113e50 .functor NAND 1, L_0x5c7c33111ce0, L_0x5c7c33111ce0, C4<1>, C4<1>;
v0x5c7c32df4500_0 .net "in_a", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df4650_0 .net "in_b", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32df4710_0 .net "out", 0 0, L_0x5c7c33113e50;  alias, 1 drivers
S_0x5c7c32df49c0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32df15b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df5100_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df51a0_0 .net "out", 0 0, L_0x5c7c33114060;  alias, 1 drivers
S_0x5c7c32df4be0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df49c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114060 .functor NAND 1, L_0x5c7c331139b0, L_0x5c7c331139b0, C4<1>, C4<1>;
v0x5c7c32df4e50_0 .net "in_a", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df4f10_0 .net "in_b", 0 0, L_0x5c7c331139b0;  alias, 1 drivers
v0x5c7c32df4fd0_0 .net "out", 0 0, L_0x5c7c33114060;  alias, 1 drivers
S_0x5c7c32df52a0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32df15b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dfad70_0 .net "branch1_out", 0 0, L_0x5c7c331143d0;  1 drivers
v0x5c7c32dfaea0_0 .net "branch2_out", 0 0, L_0x5c7c33114550;  1 drivers
v0x5c7c32dfaff0_0 .net "in_a", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
v0x5c7c32dfb0c0_0 .net "in_b", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
v0x5c7c32dfb160_0 .net "out", 0 0, L_0x5c7c331146d0;  alias, 1 drivers
v0x5c7c32dfb200_0 .net "temp1_out", 0 0, L_0x5c7c33114320;  1 drivers
v0x5c7c32dfb2a0_0 .net "temp2_out", 0 0, L_0x5c7c331144a0;  1 drivers
v0x5c7c32dfb340_0 .net "temp3_out", 0 0, L_0x5c7c33114620;  1 drivers
S_0x5c7c32df5520 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32df52a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32df65b0_0 .net "in_a", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
v0x5c7c32df6650_0 .net "in_b", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
v0x5c7c32df6710_0 .net "out", 0 0, L_0x5c7c33114320;  alias, 1 drivers
v0x5c7c32df6830_0 .net "temp_out", 0 0, L_0x5c7c33114270;  1 drivers
S_0x5c7c32df5790 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32df5520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114270 .functor NAND 1, L_0x5c7c33113fb0, L_0x5c7c33113fb0, C4<1>, C4<1>;
v0x5c7c32df5a00_0 .net "in_a", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
v0x5c7c32df5ac0_0 .net "in_b", 0 0, L_0x5c7c33113fb0;  alias, 1 drivers
v0x5c7c32df5c10_0 .net "out", 0 0, L_0x5c7c33114270;  alias, 1 drivers
S_0x5c7c32df5d10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32df5520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df6400_0 .net "in_a", 0 0, L_0x5c7c33114270;  alias, 1 drivers
v0x5c7c32df64a0_0 .net "out", 0 0, L_0x5c7c33114320;  alias, 1 drivers
S_0x5c7c32df5ee0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df5d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114320 .functor NAND 1, L_0x5c7c33114270, L_0x5c7c33114270, C4<1>, C4<1>;
v0x5c7c32df6150_0 .net "in_a", 0 0, L_0x5c7c33114270;  alias, 1 drivers
v0x5c7c32df6210_0 .net "in_b", 0 0, L_0x5c7c33114270;  alias, 1 drivers
v0x5c7c32df6300_0 .net "out", 0 0, L_0x5c7c33114320;  alias, 1 drivers
S_0x5c7c32df69a0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32df52a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32df79d0_0 .net "in_a", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
v0x5c7c32df7a70_0 .net "in_b", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
v0x5c7c32df7b30_0 .net "out", 0 0, L_0x5c7c331144a0;  alias, 1 drivers
v0x5c7c32df7c50_0 .net "temp_out", 0 0, L_0x5c7c32df97f0;  1 drivers
S_0x5c7c32df6b80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32df69a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32df97f0 .functor NAND 1, L_0x5c7c331141c0, L_0x5c7c331141c0, C4<1>, C4<1>;
v0x5c7c32df6df0_0 .net "in_a", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
v0x5c7c32df6eb0_0 .net "in_b", 0 0, L_0x5c7c331141c0;  alias, 1 drivers
v0x5c7c32df7000_0 .net "out", 0 0, L_0x5c7c32df97f0;  alias, 1 drivers
S_0x5c7c32df7100 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32df69a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df7820_0 .net "in_a", 0 0, L_0x5c7c32df97f0;  alias, 1 drivers
v0x5c7c32df78c0_0 .net "out", 0 0, L_0x5c7c331144a0;  alias, 1 drivers
S_0x5c7c32df72d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df7100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331144a0 .functor NAND 1, L_0x5c7c32df97f0, L_0x5c7c32df97f0, C4<1>, C4<1>;
v0x5c7c32df7540_0 .net "in_a", 0 0, L_0x5c7c32df97f0;  alias, 1 drivers
v0x5c7c32df7630_0 .net "in_b", 0 0, L_0x5c7c32df97f0;  alias, 1 drivers
v0x5c7c32df7720_0 .net "out", 0 0, L_0x5c7c331144a0;  alias, 1 drivers
S_0x5c7c32df7dc0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32df52a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32df8e00_0 .net "in_a", 0 0, L_0x5c7c331143d0;  alias, 1 drivers
v0x5c7c32df8ed0_0 .net "in_b", 0 0, L_0x5c7c33114550;  alias, 1 drivers
v0x5c7c32df8fa0_0 .net "out", 0 0, L_0x5c7c33114620;  alias, 1 drivers
v0x5c7c32df90c0_0 .net "temp_out", 0 0, L_0x5c7c32dfa160;  1 drivers
S_0x5c7c32df7fa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32df7dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dfa160 .functor NAND 1, L_0x5c7c331143d0, L_0x5c7c33114550, C4<1>, C4<1>;
v0x5c7c32df81f0_0 .net "in_a", 0 0, L_0x5c7c331143d0;  alias, 1 drivers
v0x5c7c32df82d0_0 .net "in_b", 0 0, L_0x5c7c33114550;  alias, 1 drivers
v0x5c7c32df8390_0 .net "out", 0 0, L_0x5c7c32dfa160;  alias, 1 drivers
S_0x5c7c32df84e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32df7dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df8c50_0 .net "in_a", 0 0, L_0x5c7c32dfa160;  alias, 1 drivers
v0x5c7c32df8cf0_0 .net "out", 0 0, L_0x5c7c33114620;  alias, 1 drivers
S_0x5c7c32df8700 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df84e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114620 .functor NAND 1, L_0x5c7c32dfa160, L_0x5c7c32dfa160, C4<1>, C4<1>;
v0x5c7c32df8970_0 .net "in_a", 0 0, L_0x5c7c32dfa160;  alias, 1 drivers
v0x5c7c32df8a60_0 .net "in_b", 0 0, L_0x5c7c32dfa160;  alias, 1 drivers
v0x5c7c32df8b50_0 .net "out", 0 0, L_0x5c7c33114620;  alias, 1 drivers
S_0x5c7c32df9210 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32df52a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32df9940_0 .net "in_a", 0 0, L_0x5c7c33114320;  alias, 1 drivers
v0x5c7c32df99e0_0 .net "out", 0 0, L_0x5c7c331143d0;  alias, 1 drivers
S_0x5c7c32df93e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df9210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331143d0 .functor NAND 1, L_0x5c7c33114320, L_0x5c7c33114320, C4<1>, C4<1>;
v0x5c7c32df9650_0 .net "in_a", 0 0, L_0x5c7c33114320;  alias, 1 drivers
v0x5c7c32df9710_0 .net "in_b", 0 0, L_0x5c7c33114320;  alias, 1 drivers
v0x5c7c32df9860_0 .net "out", 0 0, L_0x5c7c331143d0;  alias, 1 drivers
S_0x5c7c32df9ae0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32df52a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dfa2b0_0 .net "in_a", 0 0, L_0x5c7c331144a0;  alias, 1 drivers
v0x5c7c32dfa350_0 .net "out", 0 0, L_0x5c7c33114550;  alias, 1 drivers
S_0x5c7c32df9d50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32df9ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114550 .functor NAND 1, L_0x5c7c331144a0, L_0x5c7c331144a0, C4<1>, C4<1>;
v0x5c7c32df9fc0_0 .net "in_a", 0 0, L_0x5c7c331144a0;  alias, 1 drivers
v0x5c7c32dfa080_0 .net "in_b", 0 0, L_0x5c7c331144a0;  alias, 1 drivers
v0x5c7c32dfa1d0_0 .net "out", 0 0, L_0x5c7c33114550;  alias, 1 drivers
S_0x5c7c32dfa450 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32df52a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dfabf0_0 .net "in_a", 0 0, L_0x5c7c33114620;  alias, 1 drivers
v0x5c7c32dfac90_0 .net "out", 0 0, L_0x5c7c331146d0;  alias, 1 drivers
S_0x5c7c32dfa670 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dfa450;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331146d0 .functor NAND 1, L_0x5c7c33114620, L_0x5c7c33114620, C4<1>, C4<1>;
v0x5c7c32dfa8e0_0 .net "in_a", 0 0, L_0x5c7c33114620;  alias, 1 drivers
v0x5c7c32dfa9a0_0 .net "in_b", 0 0, L_0x5c7c33114620;  alias, 1 drivers
v0x5c7c32dfaaf0_0 .net "out", 0 0, L_0x5c7c331146d0;  alias, 1 drivers
S_0x5c7c32dfbef0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32de3d30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e018e0_0 .net "branch1_out", 0 0, L_0x5c7c33114960;  1 drivers
v0x5c7c32e01a10_0 .net "branch2_out", 0 0, L_0x5c7c33114bf0;  1 drivers
v0x5c7c32e01b60_0 .net "in_a", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32e01d40_0 .net "in_b", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32e01ef0_0 .net "out", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e01f90_0 .net "temp1_out", 0 0, L_0x5c7c331148b0;  1 drivers
v0x5c7c32e02030_0 .net "temp2_out", 0 0, L_0x5c7c33114b40;  1 drivers
v0x5c7c32e020d0_0 .net "temp3_out", 0 0, L_0x5c7c33114dd0;  1 drivers
S_0x5c7c32dfc080 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32dfbef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dfd120_0 .net "in_a", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32dfd1c0_0 .net "in_b", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32dfd280_0 .net "out", 0 0, L_0x5c7c331148b0;  alias, 1 drivers
v0x5c7c32dfd3a0_0 .net "temp_out", 0 0, L_0x5c7c32dfaa80;  1 drivers
S_0x5c7c32dfc2a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dfc080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32dfaa80 .functor NAND 1, L_0x5c7c33112d40, L_0x5c7c33112d40, C4<1>, C4<1>;
v0x5c7c32dfc510_0 .net "in_a", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32dfc660_0 .net "in_b", 0 0, L_0x5c7c33112d40;  alias, 1 drivers
v0x5c7c32dfc720_0 .net "out", 0 0, L_0x5c7c32dfaa80;  alias, 1 drivers
S_0x5c7c32dfc850 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dfc080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dfcf70_0 .net "in_a", 0 0, L_0x5c7c32dfaa80;  alias, 1 drivers
v0x5c7c32dfd010_0 .net "out", 0 0, L_0x5c7c331148b0;  alias, 1 drivers
S_0x5c7c32dfca20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dfc850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331148b0 .functor NAND 1, L_0x5c7c32dfaa80, L_0x5c7c32dfaa80, C4<1>, C4<1>;
v0x5c7c32dfcc90_0 .net "in_a", 0 0, L_0x5c7c32dfaa80;  alias, 1 drivers
v0x5c7c32dfcd80_0 .net "in_b", 0 0, L_0x5c7c32dfaa80;  alias, 1 drivers
v0x5c7c32dfce70_0 .net "out", 0 0, L_0x5c7c331148b0;  alias, 1 drivers
S_0x5c7c32dfd510 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32dfbef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dfe540_0 .net "in_a", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32dfe5e0_0 .net "in_b", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32dfe6a0_0 .net "out", 0 0, L_0x5c7c33114b40;  alias, 1 drivers
v0x5c7c32dfe7c0_0 .net "temp_out", 0 0, L_0x5c7c32e00360;  1 drivers
S_0x5c7c32dfd6f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dfd510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e00360 .functor NAND 1, L_0x5c7c33113da0, L_0x5c7c33113da0, C4<1>, C4<1>;
v0x5c7c32dfd960_0 .net "in_a", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32dfdab0_0 .net "in_b", 0 0, L_0x5c7c33113da0;  alias, 1 drivers
v0x5c7c32dfdb70_0 .net "out", 0 0, L_0x5c7c32e00360;  alias, 1 drivers
S_0x5c7c32dfdc70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dfd510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dfe390_0 .net "in_a", 0 0, L_0x5c7c32e00360;  alias, 1 drivers
v0x5c7c32dfe430_0 .net "out", 0 0, L_0x5c7c33114b40;  alias, 1 drivers
S_0x5c7c32dfde40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dfdc70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114b40 .functor NAND 1, L_0x5c7c32e00360, L_0x5c7c32e00360, C4<1>, C4<1>;
v0x5c7c32dfe0b0_0 .net "in_a", 0 0, L_0x5c7c32e00360;  alias, 1 drivers
v0x5c7c32dfe1a0_0 .net "in_b", 0 0, L_0x5c7c32e00360;  alias, 1 drivers
v0x5c7c32dfe290_0 .net "out", 0 0, L_0x5c7c33114b40;  alias, 1 drivers
S_0x5c7c32dfe930 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32dfbef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32dff970_0 .net "in_a", 0 0, L_0x5c7c33114960;  alias, 1 drivers
v0x5c7c32dffa40_0 .net "in_b", 0 0, L_0x5c7c33114bf0;  alias, 1 drivers
v0x5c7c32dffb10_0 .net "out", 0 0, L_0x5c7c33114dd0;  alias, 1 drivers
v0x5c7c32dffc30_0 .net "temp_out", 0 0, L_0x5c7c32e00cd0;  1 drivers
S_0x5c7c32dfeb10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32dfe930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e00cd0 .functor NAND 1, L_0x5c7c33114960, L_0x5c7c33114bf0, C4<1>, C4<1>;
v0x5c7c32dfed60_0 .net "in_a", 0 0, L_0x5c7c33114960;  alias, 1 drivers
v0x5c7c32dfee40_0 .net "in_b", 0 0, L_0x5c7c33114bf0;  alias, 1 drivers
v0x5c7c32dfef00_0 .net "out", 0 0, L_0x5c7c32e00cd0;  alias, 1 drivers
S_0x5c7c32dff050 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32dfe930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32dff7c0_0 .net "in_a", 0 0, L_0x5c7c32e00cd0;  alias, 1 drivers
v0x5c7c32dff860_0 .net "out", 0 0, L_0x5c7c33114dd0;  alias, 1 drivers
S_0x5c7c32dff270 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dff050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114dd0 .functor NAND 1, L_0x5c7c32e00cd0, L_0x5c7c32e00cd0, C4<1>, C4<1>;
v0x5c7c32dff4e0_0 .net "in_a", 0 0, L_0x5c7c32e00cd0;  alias, 1 drivers
v0x5c7c32dff5d0_0 .net "in_b", 0 0, L_0x5c7c32e00cd0;  alias, 1 drivers
v0x5c7c32dff6c0_0 .net "out", 0 0, L_0x5c7c33114dd0;  alias, 1 drivers
S_0x5c7c32dffd80 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32dfbef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e004b0_0 .net "in_a", 0 0, L_0x5c7c331148b0;  alias, 1 drivers
v0x5c7c32e00550_0 .net "out", 0 0, L_0x5c7c33114960;  alias, 1 drivers
S_0x5c7c32dfff50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32dffd80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114960 .functor NAND 1, L_0x5c7c331148b0, L_0x5c7c331148b0, C4<1>, C4<1>;
v0x5c7c32e001c0_0 .net "in_a", 0 0, L_0x5c7c331148b0;  alias, 1 drivers
v0x5c7c32e00280_0 .net "in_b", 0 0, L_0x5c7c331148b0;  alias, 1 drivers
v0x5c7c32e003d0_0 .net "out", 0 0, L_0x5c7c33114960;  alias, 1 drivers
S_0x5c7c32e00650 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32dfbef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e00e20_0 .net "in_a", 0 0, L_0x5c7c33114b40;  alias, 1 drivers
v0x5c7c32e00ec0_0 .net "out", 0 0, L_0x5c7c33114bf0;  alias, 1 drivers
S_0x5c7c32e008c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e00650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114bf0 .functor NAND 1, L_0x5c7c33114b40, L_0x5c7c33114b40, C4<1>, C4<1>;
v0x5c7c32e00b30_0 .net "in_a", 0 0, L_0x5c7c33114b40;  alias, 1 drivers
v0x5c7c32e00bf0_0 .net "in_b", 0 0, L_0x5c7c33114b40;  alias, 1 drivers
v0x5c7c32e00d40_0 .net "out", 0 0, L_0x5c7c33114bf0;  alias, 1 drivers
S_0x5c7c32e00fc0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32dfbef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e01760_0 .net "in_a", 0 0, L_0x5c7c33114dd0;  alias, 1 drivers
v0x5c7c32e01800_0 .net "out", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
S_0x5c7c32e011e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e00fc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33114e80 .functor NAND 1, L_0x5c7c33114dd0, L_0x5c7c33114dd0, C4<1>, C4<1>;
v0x5c7c32e01450_0 .net "in_a", 0 0, L_0x5c7c33114dd0;  alias, 1 drivers
v0x5c7c32e01510_0 .net "in_b", 0 0, L_0x5c7c33114dd0;  alias, 1 drivers
v0x5c7c32e01660_0 .net "out", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
S_0x5c7c32e02730 .scope module, "fa_gate3" "FullAdder" 2 8, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32e20ba0_0 .net "a", 0 0, L_0x5c7c33117620;  1 drivers
v0x5c7c32e20c40_0 .net "b", 0 0, L_0x5c7c331176c0;  1 drivers
v0x5c7c32e20d00_0 .net "c", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e20da0_0 .net "carry", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e20e40_0 .net "sum", 0 0, L_0x5c7c33116cd0;  1 drivers
v0x5c7c32e20ee0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33115250;  1 drivers
v0x5c7c32e20f80_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c331163a0;  1 drivers
v0x5c7c32e21020_0 .net "tmp_sum_out", 0 0, L_0x5c7c33115da0;  1 drivers
S_0x5c7c32e02990 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32e02730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e0e550_0 .net "a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e0e700_0 .net "b", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e0e8d0_0 .net "carry", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e0e970_0 .net "sum", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
S_0x5c7c32e02bb0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e02990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e03ca0_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e03d70_0 .net "in_b", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e03e40_0 .net "out", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e03f60_0 .net "temp_out", 0 0, L_0x5c7c331151e0;  1 drivers
S_0x5c7c32e02e20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e02bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331151e0 .functor NAND 1, L_0x5c7c33117620, L_0x5c7c331176c0, C4<1>, C4<1>;
v0x5c7c32e03090_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e03170_0 .net "in_b", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e03230_0 .net "out", 0 0, L_0x5c7c331151e0;  alias, 1 drivers
S_0x5c7c32e03380 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e02bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e03af0_0 .net "in_a", 0 0, L_0x5c7c331151e0;  alias, 1 drivers
v0x5c7c32e03b90_0 .net "out", 0 0, L_0x5c7c33115250;  alias, 1 drivers
S_0x5c7c32e035a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e03380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115250 .functor NAND 1, L_0x5c7c331151e0, L_0x5c7c331151e0, C4<1>, C4<1>;
v0x5c7c32e03810_0 .net "in_a", 0 0, L_0x5c7c331151e0;  alias, 1 drivers
v0x5c7c32e03900_0 .net "in_b", 0 0, L_0x5c7c331151e0;  alias, 1 drivers
v0x5c7c32e039f0_0 .net "out", 0 0, L_0x5c7c33115250;  alias, 1 drivers
S_0x5c7c32e04020 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e02990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e0de70_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e0df10_0 .net "in_b", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e0dfd0_0 .net "out", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e0e070_0 .net "temp_a_and_out", 0 0, L_0x5c7c33115460;  1 drivers
v0x5c7c32e0e220_0 .net "temp_a_out", 0 0, L_0x5c7c33115300;  1 drivers
v0x5c7c32e0e2c0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33115670;  1 drivers
v0x5c7c32e0e470_0 .net "temp_b_out", 0 0, L_0x5c7c33115510;  1 drivers
S_0x5c7c32e04200 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e04020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e052c0_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e05360_0 .net "in_b", 0 0, L_0x5c7c33115300;  alias, 1 drivers
v0x5c7c32e05450_0 .net "out", 0 0, L_0x5c7c33115460;  alias, 1 drivers
v0x5c7c32e05570_0 .net "temp_out", 0 0, L_0x5c7c331153b0;  1 drivers
S_0x5c7c32e04470 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e04200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331153b0 .functor NAND 1, L_0x5c7c33117620, L_0x5c7c33115300, C4<1>, C4<1>;
v0x5c7c32e046e0_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e047f0_0 .net "in_b", 0 0, L_0x5c7c33115300;  alias, 1 drivers
v0x5c7c32e048b0_0 .net "out", 0 0, L_0x5c7c331153b0;  alias, 1 drivers
S_0x5c7c32e049d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e04200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e05110_0 .net "in_a", 0 0, L_0x5c7c331153b0;  alias, 1 drivers
v0x5c7c32e051b0_0 .net "out", 0 0, L_0x5c7c33115460;  alias, 1 drivers
S_0x5c7c32e04bf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e049d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115460 .functor NAND 1, L_0x5c7c331153b0, L_0x5c7c331153b0, C4<1>, C4<1>;
v0x5c7c32e04e60_0 .net "in_a", 0 0, L_0x5c7c331153b0;  alias, 1 drivers
v0x5c7c32e04f20_0 .net "in_b", 0 0, L_0x5c7c331153b0;  alias, 1 drivers
v0x5c7c32e05010_0 .net "out", 0 0, L_0x5c7c33115460;  alias, 1 drivers
S_0x5c7c32e056c0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e04020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e066f0_0 .net "in_a", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e06790_0 .net "in_b", 0 0, L_0x5c7c33115510;  alias, 1 drivers
v0x5c7c32e06880_0 .net "out", 0 0, L_0x5c7c33115670;  alias, 1 drivers
v0x5c7c32e069a0_0 .net "temp_out", 0 0, L_0x5c7c331155c0;  1 drivers
S_0x5c7c32e058a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e056c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331155c0 .functor NAND 1, L_0x5c7c331176c0, L_0x5c7c33115510, C4<1>, C4<1>;
v0x5c7c32e05b10_0 .net "in_a", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e05c20_0 .net "in_b", 0 0, L_0x5c7c33115510;  alias, 1 drivers
v0x5c7c32e05ce0_0 .net "out", 0 0, L_0x5c7c331155c0;  alias, 1 drivers
S_0x5c7c32e05e00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e056c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e06540_0 .net "in_a", 0 0, L_0x5c7c331155c0;  alias, 1 drivers
v0x5c7c32e065e0_0 .net "out", 0 0, L_0x5c7c33115670;  alias, 1 drivers
S_0x5c7c32e06020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e05e00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115670 .functor NAND 1, L_0x5c7c331155c0, L_0x5c7c331155c0, C4<1>, C4<1>;
v0x5c7c32e06290_0 .net "in_a", 0 0, L_0x5c7c331155c0;  alias, 1 drivers
v0x5c7c32e06350_0 .net "in_b", 0 0, L_0x5c7c331155c0;  alias, 1 drivers
v0x5c7c32e06440_0 .net "out", 0 0, L_0x5c7c33115670;  alias, 1 drivers
S_0x5c7c32e06af0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e04020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e07230_0 .net "in_a", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e072d0_0 .net "out", 0 0, L_0x5c7c33115300;  alias, 1 drivers
S_0x5c7c32e06cc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e06af0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115300 .functor NAND 1, L_0x5c7c331176c0, L_0x5c7c331176c0, C4<1>, C4<1>;
v0x5c7c32e06f10_0 .net "in_a", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e07060_0 .net "in_b", 0 0, L_0x5c7c331176c0;  alias, 1 drivers
v0x5c7c32e07120_0 .net "out", 0 0, L_0x5c7c33115300;  alias, 1 drivers
S_0x5c7c32e073d0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e04020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e07b50_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e07bf0_0 .net "out", 0 0, L_0x5c7c33115510;  alias, 1 drivers
S_0x5c7c32e075f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e073d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115510 .functor NAND 1, L_0x5c7c33117620, L_0x5c7c33117620, C4<1>, C4<1>;
v0x5c7c32e07860_0 .net "in_a", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e079b0_0 .net "in_b", 0 0, L_0x5c7c33117620;  alias, 1 drivers
v0x5c7c32e07a70_0 .net "out", 0 0, L_0x5c7c33115510;  alias, 1 drivers
S_0x5c7c32e07cf0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e04020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e0d7c0_0 .net "branch1_out", 0 0, L_0x5c7c33115880;  1 drivers
v0x5c7c32e0d8f0_0 .net "branch2_out", 0 0, L_0x5c7c33115b10;  1 drivers
v0x5c7c32e0da40_0 .net "in_a", 0 0, L_0x5c7c33115460;  alias, 1 drivers
v0x5c7c32e0db10_0 .net "in_b", 0 0, L_0x5c7c33115670;  alias, 1 drivers
v0x5c7c32e0dbb0_0 .net "out", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e0dc50_0 .net "temp1_out", 0 0, L_0x5c7c331157d0;  1 drivers
v0x5c7c32e0dcf0_0 .net "temp2_out", 0 0, L_0x5c7c33115a60;  1 drivers
v0x5c7c32e0dd90_0 .net "temp3_out", 0 0, L_0x5c7c33115cf0;  1 drivers
S_0x5c7c32e07f70 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e07cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e09000_0 .net "in_a", 0 0, L_0x5c7c33115460;  alias, 1 drivers
v0x5c7c32e090a0_0 .net "in_b", 0 0, L_0x5c7c33115460;  alias, 1 drivers
v0x5c7c32e09160_0 .net "out", 0 0, L_0x5c7c331157d0;  alias, 1 drivers
v0x5c7c32e09280_0 .net "temp_out", 0 0, L_0x5c7c33115720;  1 drivers
S_0x5c7c32e081e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e07f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115720 .functor NAND 1, L_0x5c7c33115460, L_0x5c7c33115460, C4<1>, C4<1>;
v0x5c7c32e08450_0 .net "in_a", 0 0, L_0x5c7c33115460;  alias, 1 drivers
v0x5c7c32e08510_0 .net "in_b", 0 0, L_0x5c7c33115460;  alias, 1 drivers
v0x5c7c32e08660_0 .net "out", 0 0, L_0x5c7c33115720;  alias, 1 drivers
S_0x5c7c32e08760 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e07f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e08e50_0 .net "in_a", 0 0, L_0x5c7c33115720;  alias, 1 drivers
v0x5c7c32e08ef0_0 .net "out", 0 0, L_0x5c7c331157d0;  alias, 1 drivers
S_0x5c7c32e08930 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e08760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331157d0 .functor NAND 1, L_0x5c7c33115720, L_0x5c7c33115720, C4<1>, C4<1>;
v0x5c7c32e08ba0_0 .net "in_a", 0 0, L_0x5c7c33115720;  alias, 1 drivers
v0x5c7c32e08c60_0 .net "in_b", 0 0, L_0x5c7c33115720;  alias, 1 drivers
v0x5c7c32e08d50_0 .net "out", 0 0, L_0x5c7c331157d0;  alias, 1 drivers
S_0x5c7c32e093f0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e07cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e0a420_0 .net "in_a", 0 0, L_0x5c7c33115670;  alias, 1 drivers
v0x5c7c32e0a4c0_0 .net "in_b", 0 0, L_0x5c7c33115670;  alias, 1 drivers
v0x5c7c32e0a580_0 .net "out", 0 0, L_0x5c7c33115a60;  alias, 1 drivers
v0x5c7c32e0a6a0_0 .net "temp_out", 0 0, L_0x5c7c32e0c240;  1 drivers
S_0x5c7c32e095d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e093f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e0c240 .functor NAND 1, L_0x5c7c33115670, L_0x5c7c33115670, C4<1>, C4<1>;
v0x5c7c32e09840_0 .net "in_a", 0 0, L_0x5c7c33115670;  alias, 1 drivers
v0x5c7c32e09900_0 .net "in_b", 0 0, L_0x5c7c33115670;  alias, 1 drivers
v0x5c7c32e09a50_0 .net "out", 0 0, L_0x5c7c32e0c240;  alias, 1 drivers
S_0x5c7c32e09b50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e093f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e0a270_0 .net "in_a", 0 0, L_0x5c7c32e0c240;  alias, 1 drivers
v0x5c7c32e0a310_0 .net "out", 0 0, L_0x5c7c33115a60;  alias, 1 drivers
S_0x5c7c32e09d20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e09b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115a60 .functor NAND 1, L_0x5c7c32e0c240, L_0x5c7c32e0c240, C4<1>, C4<1>;
v0x5c7c32e09f90_0 .net "in_a", 0 0, L_0x5c7c32e0c240;  alias, 1 drivers
v0x5c7c32e0a080_0 .net "in_b", 0 0, L_0x5c7c32e0c240;  alias, 1 drivers
v0x5c7c32e0a170_0 .net "out", 0 0, L_0x5c7c33115a60;  alias, 1 drivers
S_0x5c7c32e0a810 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e07cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e0b850_0 .net "in_a", 0 0, L_0x5c7c33115880;  alias, 1 drivers
v0x5c7c32e0b920_0 .net "in_b", 0 0, L_0x5c7c33115b10;  alias, 1 drivers
v0x5c7c32e0b9f0_0 .net "out", 0 0, L_0x5c7c33115cf0;  alias, 1 drivers
v0x5c7c32e0bb10_0 .net "temp_out", 0 0, L_0x5c7c32e0cbb0;  1 drivers
S_0x5c7c32e0a9f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e0a810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e0cbb0 .functor NAND 1, L_0x5c7c33115880, L_0x5c7c33115b10, C4<1>, C4<1>;
v0x5c7c32e0ac40_0 .net "in_a", 0 0, L_0x5c7c33115880;  alias, 1 drivers
v0x5c7c32e0ad20_0 .net "in_b", 0 0, L_0x5c7c33115b10;  alias, 1 drivers
v0x5c7c32e0ade0_0 .net "out", 0 0, L_0x5c7c32e0cbb0;  alias, 1 drivers
S_0x5c7c32e0af30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e0a810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e0b6a0_0 .net "in_a", 0 0, L_0x5c7c32e0cbb0;  alias, 1 drivers
v0x5c7c32e0b740_0 .net "out", 0 0, L_0x5c7c33115cf0;  alias, 1 drivers
S_0x5c7c32e0b150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e0af30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115cf0 .functor NAND 1, L_0x5c7c32e0cbb0, L_0x5c7c32e0cbb0, C4<1>, C4<1>;
v0x5c7c32e0b3c0_0 .net "in_a", 0 0, L_0x5c7c32e0cbb0;  alias, 1 drivers
v0x5c7c32e0b4b0_0 .net "in_b", 0 0, L_0x5c7c32e0cbb0;  alias, 1 drivers
v0x5c7c32e0b5a0_0 .net "out", 0 0, L_0x5c7c33115cf0;  alias, 1 drivers
S_0x5c7c32e0bc60 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e07cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e0c390_0 .net "in_a", 0 0, L_0x5c7c331157d0;  alias, 1 drivers
v0x5c7c32e0c430_0 .net "out", 0 0, L_0x5c7c33115880;  alias, 1 drivers
S_0x5c7c32e0be30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e0bc60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115880 .functor NAND 1, L_0x5c7c331157d0, L_0x5c7c331157d0, C4<1>, C4<1>;
v0x5c7c32e0c0a0_0 .net "in_a", 0 0, L_0x5c7c331157d0;  alias, 1 drivers
v0x5c7c32e0c160_0 .net "in_b", 0 0, L_0x5c7c331157d0;  alias, 1 drivers
v0x5c7c32e0c2b0_0 .net "out", 0 0, L_0x5c7c33115880;  alias, 1 drivers
S_0x5c7c32e0c530 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e07cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e0cd00_0 .net "in_a", 0 0, L_0x5c7c33115a60;  alias, 1 drivers
v0x5c7c32e0cda0_0 .net "out", 0 0, L_0x5c7c33115b10;  alias, 1 drivers
S_0x5c7c32e0c7a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e0c530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115b10 .functor NAND 1, L_0x5c7c33115a60, L_0x5c7c33115a60, C4<1>, C4<1>;
v0x5c7c32e0ca10_0 .net "in_a", 0 0, L_0x5c7c33115a60;  alias, 1 drivers
v0x5c7c32e0cad0_0 .net "in_b", 0 0, L_0x5c7c33115a60;  alias, 1 drivers
v0x5c7c32e0cc20_0 .net "out", 0 0, L_0x5c7c33115b10;  alias, 1 drivers
S_0x5c7c32e0cea0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e07cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e0d640_0 .net "in_a", 0 0, L_0x5c7c33115cf0;  alias, 1 drivers
v0x5c7c32e0d6e0_0 .net "out", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
S_0x5c7c32e0d0c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e0cea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33115da0 .functor NAND 1, L_0x5c7c33115cf0, L_0x5c7c33115cf0, C4<1>, C4<1>;
v0x5c7c32e0d330_0 .net "in_a", 0 0, L_0x5c7c33115cf0;  alias, 1 drivers
v0x5c7c32e0d3f0_0 .net "in_b", 0 0, L_0x5c7c33115cf0;  alias, 1 drivers
v0x5c7c32e0d540_0 .net "out", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
S_0x5c7c32e0ea50 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32e02730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e1a570_0 .net "a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e1a610_0 .net "b", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e1a6d0_0 .net "carry", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e1a770_0 .net "sum", 0 0, L_0x5c7c33116cd0;  alias, 1 drivers
S_0x5c7c32e0ec70 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e0ea50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e0fc10_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e0fcb0_0 .net "in_b", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e0fd70_0 .net "out", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e0fe90_0 .net "temp_out", 0 0, L_0x5c7c32e0d4d0;  1 drivers
S_0x5c7c32e0ee20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e0ec70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e0d4d0 .functor NAND 1, L_0x5c7c33115da0, L_0x5c7c33114e80, C4<1>, C4<1>;
v0x5c7c32e0f090_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e0f150_0 .net "in_b", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e0f210_0 .net "out", 0 0, L_0x5c7c32e0d4d0;  alias, 1 drivers
S_0x5c7c32e0f340 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e0ec70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e0fa60_0 .net "in_a", 0 0, L_0x5c7c32e0d4d0;  alias, 1 drivers
v0x5c7c32e0fb00_0 .net "out", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
S_0x5c7c32e0f510 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e0f340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331163a0 .functor NAND 1, L_0x5c7c32e0d4d0, L_0x5c7c32e0d4d0, C4<1>, C4<1>;
v0x5c7c32e0f780_0 .net "in_a", 0 0, L_0x5c7c32e0d4d0;  alias, 1 drivers
v0x5c7c32e0f870_0 .net "in_b", 0 0, L_0x5c7c32e0d4d0;  alias, 1 drivers
v0x5c7c32e0f960_0 .net "out", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
S_0x5c7c32e10000 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e0ea50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e19e90_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e19f30_0 .net "in_b", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e19ff0_0 .net "out", 0 0, L_0x5c7c33116cd0;  alias, 1 drivers
v0x5c7c32e1a090_0 .net "temp_a_and_out", 0 0, L_0x5c7c331165b0;  1 drivers
v0x5c7c32e1a240_0 .net "temp_a_out", 0 0, L_0x5c7c33116450;  1 drivers
v0x5c7c32e1a2e0_0 .net "temp_b_and_out", 0 0, L_0x5c7c331167c0;  1 drivers
v0x5c7c32e1a490_0 .net "temp_b_out", 0 0, L_0x5c7c33116660;  1 drivers
S_0x5c7c32e101e0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e10000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e11280_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e11430_0 .net "in_b", 0 0, L_0x5c7c33116450;  alias, 1 drivers
v0x5c7c32e11520_0 .net "out", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
v0x5c7c32e11640_0 .net "temp_out", 0 0, L_0x5c7c33116500;  1 drivers
S_0x5c7c32e10450 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e101e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116500 .functor NAND 1, L_0x5c7c33115da0, L_0x5c7c33116450, C4<1>, C4<1>;
v0x5c7c32e106c0_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e10780_0 .net "in_b", 0 0, L_0x5c7c33116450;  alias, 1 drivers
v0x5c7c32e10840_0 .net "out", 0 0, L_0x5c7c33116500;  alias, 1 drivers
S_0x5c7c32e10960 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e101e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e110d0_0 .net "in_a", 0 0, L_0x5c7c33116500;  alias, 1 drivers
v0x5c7c32e11170_0 .net "out", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
S_0x5c7c32e10b80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e10960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331165b0 .functor NAND 1, L_0x5c7c33116500, L_0x5c7c33116500, C4<1>, C4<1>;
v0x5c7c32e10df0_0 .net "in_a", 0 0, L_0x5c7c33116500;  alias, 1 drivers
v0x5c7c32e10ee0_0 .net "in_b", 0 0, L_0x5c7c33116500;  alias, 1 drivers
v0x5c7c32e10fd0_0 .net "out", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
S_0x5c7c32e11700 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e10000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e12710_0 .net "in_a", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e127b0_0 .net "in_b", 0 0, L_0x5c7c33116660;  alias, 1 drivers
v0x5c7c32e128a0_0 .net "out", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
v0x5c7c32e129c0_0 .net "temp_out", 0 0, L_0x5c7c33116710;  1 drivers
S_0x5c7c32e118e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e11700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116710 .functor NAND 1, L_0x5c7c33114e80, L_0x5c7c33116660, C4<1>, C4<1>;
v0x5c7c32e11b50_0 .net "in_a", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e11c10_0 .net "in_b", 0 0, L_0x5c7c33116660;  alias, 1 drivers
v0x5c7c32e11cd0_0 .net "out", 0 0, L_0x5c7c33116710;  alias, 1 drivers
S_0x5c7c32e11df0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e11700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e12560_0 .net "in_a", 0 0, L_0x5c7c33116710;  alias, 1 drivers
v0x5c7c32e12600_0 .net "out", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
S_0x5c7c32e12010 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e11df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331167c0 .functor NAND 1, L_0x5c7c33116710, L_0x5c7c33116710, C4<1>, C4<1>;
v0x5c7c32e12280_0 .net "in_a", 0 0, L_0x5c7c33116710;  alias, 1 drivers
v0x5c7c32e12370_0 .net "in_b", 0 0, L_0x5c7c33116710;  alias, 1 drivers
v0x5c7c32e12460_0 .net "out", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
S_0x5c7c32e12b10 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e10000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e13320_0 .net "in_a", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e133c0_0 .net "out", 0 0, L_0x5c7c33116450;  alias, 1 drivers
S_0x5c7c32e12ce0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e12b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116450 .functor NAND 1, L_0x5c7c33114e80, L_0x5c7c33114e80, C4<1>, C4<1>;
v0x5c7c32e12f30_0 .net "in_a", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e13100_0 .net "in_b", 0 0, L_0x5c7c33114e80;  alias, 1 drivers
v0x5c7c32e131c0_0 .net "out", 0 0, L_0x5c7c33116450;  alias, 1 drivers
S_0x5c7c32e134c0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e10000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e13c00_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e13ca0_0 .net "out", 0 0, L_0x5c7c33116660;  alias, 1 drivers
S_0x5c7c32e136e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e134c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116660 .functor NAND 1, L_0x5c7c33115da0, L_0x5c7c33115da0, C4<1>, C4<1>;
v0x5c7c32e13950_0 .net "in_a", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e13a10_0 .net "in_b", 0 0, L_0x5c7c33115da0;  alias, 1 drivers
v0x5c7c32e13ad0_0 .net "out", 0 0, L_0x5c7c33116660;  alias, 1 drivers
S_0x5c7c32e13da0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e10000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e197e0_0 .net "branch1_out", 0 0, L_0x5c7c331169d0;  1 drivers
v0x5c7c32e19910_0 .net "branch2_out", 0 0, L_0x5c7c33116b50;  1 drivers
v0x5c7c32e19a60_0 .net "in_a", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
v0x5c7c32e19b30_0 .net "in_b", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
v0x5c7c32e19bd0_0 .net "out", 0 0, L_0x5c7c33116cd0;  alias, 1 drivers
v0x5c7c32e19c70_0 .net "temp1_out", 0 0, L_0x5c7c33116920;  1 drivers
v0x5c7c32e19d10_0 .net "temp2_out", 0 0, L_0x5c7c33116aa0;  1 drivers
v0x5c7c32e19db0_0 .net "temp3_out", 0 0, L_0x5c7c33116c20;  1 drivers
S_0x5c7c32e14020 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e13da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e15020_0 .net "in_a", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
v0x5c7c32e150c0_0 .net "in_b", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
v0x5c7c32e15180_0 .net "out", 0 0, L_0x5c7c33116920;  alias, 1 drivers
v0x5c7c32e152a0_0 .net "temp_out", 0 0, L_0x5c7c33116870;  1 drivers
S_0x5c7c32e14290 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e14020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116870 .functor NAND 1, L_0x5c7c331165b0, L_0x5c7c331165b0, C4<1>, C4<1>;
v0x5c7c32e14500_0 .net "in_a", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
v0x5c7c32e145c0_0 .net "in_b", 0 0, L_0x5c7c331165b0;  alias, 1 drivers
v0x5c7c32e14680_0 .net "out", 0 0, L_0x5c7c33116870;  alias, 1 drivers
S_0x5c7c32e14780 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e14020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e14e70_0 .net "in_a", 0 0, L_0x5c7c33116870;  alias, 1 drivers
v0x5c7c32e14f10_0 .net "out", 0 0, L_0x5c7c33116920;  alias, 1 drivers
S_0x5c7c32e14950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e14780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116920 .functor NAND 1, L_0x5c7c33116870, L_0x5c7c33116870, C4<1>, C4<1>;
v0x5c7c32e14bc0_0 .net "in_a", 0 0, L_0x5c7c33116870;  alias, 1 drivers
v0x5c7c32e14c80_0 .net "in_b", 0 0, L_0x5c7c33116870;  alias, 1 drivers
v0x5c7c32e14d70_0 .net "out", 0 0, L_0x5c7c33116920;  alias, 1 drivers
S_0x5c7c32e15410 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e13da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e16440_0 .net "in_a", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
v0x5c7c32e164e0_0 .net "in_b", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
v0x5c7c32e165a0_0 .net "out", 0 0, L_0x5c7c33116aa0;  alias, 1 drivers
v0x5c7c32e166c0_0 .net "temp_out", 0 0, L_0x5c7c32e18260;  1 drivers
S_0x5c7c32e155f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e15410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e18260 .functor NAND 1, L_0x5c7c331167c0, L_0x5c7c331167c0, C4<1>, C4<1>;
v0x5c7c32e15860_0 .net "in_a", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
v0x5c7c32e15920_0 .net "in_b", 0 0, L_0x5c7c331167c0;  alias, 1 drivers
v0x5c7c32e15a70_0 .net "out", 0 0, L_0x5c7c32e18260;  alias, 1 drivers
S_0x5c7c32e15b70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e15410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e16290_0 .net "in_a", 0 0, L_0x5c7c32e18260;  alias, 1 drivers
v0x5c7c32e16330_0 .net "out", 0 0, L_0x5c7c33116aa0;  alias, 1 drivers
S_0x5c7c32e15d40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e15b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116aa0 .functor NAND 1, L_0x5c7c32e18260, L_0x5c7c32e18260, C4<1>, C4<1>;
v0x5c7c32e15fb0_0 .net "in_a", 0 0, L_0x5c7c32e18260;  alias, 1 drivers
v0x5c7c32e160a0_0 .net "in_b", 0 0, L_0x5c7c32e18260;  alias, 1 drivers
v0x5c7c32e16190_0 .net "out", 0 0, L_0x5c7c33116aa0;  alias, 1 drivers
S_0x5c7c32e16830 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e13da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e17870_0 .net "in_a", 0 0, L_0x5c7c331169d0;  alias, 1 drivers
v0x5c7c32e17940_0 .net "in_b", 0 0, L_0x5c7c33116b50;  alias, 1 drivers
v0x5c7c32e17a10_0 .net "out", 0 0, L_0x5c7c33116c20;  alias, 1 drivers
v0x5c7c32e17b30_0 .net "temp_out", 0 0, L_0x5c7c32e18bd0;  1 drivers
S_0x5c7c32e16a10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e16830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e18bd0 .functor NAND 1, L_0x5c7c331169d0, L_0x5c7c33116b50, C4<1>, C4<1>;
v0x5c7c32e16c60_0 .net "in_a", 0 0, L_0x5c7c331169d0;  alias, 1 drivers
v0x5c7c32e16d40_0 .net "in_b", 0 0, L_0x5c7c33116b50;  alias, 1 drivers
v0x5c7c32e16e00_0 .net "out", 0 0, L_0x5c7c32e18bd0;  alias, 1 drivers
S_0x5c7c32e16f50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e16830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e176c0_0 .net "in_a", 0 0, L_0x5c7c32e18bd0;  alias, 1 drivers
v0x5c7c32e17760_0 .net "out", 0 0, L_0x5c7c33116c20;  alias, 1 drivers
S_0x5c7c32e17170 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e16f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116c20 .functor NAND 1, L_0x5c7c32e18bd0, L_0x5c7c32e18bd0, C4<1>, C4<1>;
v0x5c7c32e173e0_0 .net "in_a", 0 0, L_0x5c7c32e18bd0;  alias, 1 drivers
v0x5c7c32e174d0_0 .net "in_b", 0 0, L_0x5c7c32e18bd0;  alias, 1 drivers
v0x5c7c32e175c0_0 .net "out", 0 0, L_0x5c7c33116c20;  alias, 1 drivers
S_0x5c7c32e17c80 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e13da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e183b0_0 .net "in_a", 0 0, L_0x5c7c33116920;  alias, 1 drivers
v0x5c7c32e18450_0 .net "out", 0 0, L_0x5c7c331169d0;  alias, 1 drivers
S_0x5c7c32e17e50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e17c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331169d0 .functor NAND 1, L_0x5c7c33116920, L_0x5c7c33116920, C4<1>, C4<1>;
v0x5c7c32e180c0_0 .net "in_a", 0 0, L_0x5c7c33116920;  alias, 1 drivers
v0x5c7c32e18180_0 .net "in_b", 0 0, L_0x5c7c33116920;  alias, 1 drivers
v0x5c7c32e182d0_0 .net "out", 0 0, L_0x5c7c331169d0;  alias, 1 drivers
S_0x5c7c32e18550 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e13da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e18d20_0 .net "in_a", 0 0, L_0x5c7c33116aa0;  alias, 1 drivers
v0x5c7c32e18dc0_0 .net "out", 0 0, L_0x5c7c33116b50;  alias, 1 drivers
S_0x5c7c32e187c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e18550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116b50 .functor NAND 1, L_0x5c7c33116aa0, L_0x5c7c33116aa0, C4<1>, C4<1>;
v0x5c7c32e18a30_0 .net "in_a", 0 0, L_0x5c7c33116aa0;  alias, 1 drivers
v0x5c7c32e18af0_0 .net "in_b", 0 0, L_0x5c7c33116aa0;  alias, 1 drivers
v0x5c7c32e18c40_0 .net "out", 0 0, L_0x5c7c33116b50;  alias, 1 drivers
S_0x5c7c32e18ec0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e13da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e19660_0 .net "in_a", 0 0, L_0x5c7c33116c20;  alias, 1 drivers
v0x5c7c32e19700_0 .net "out", 0 0, L_0x5c7c33116cd0;  alias, 1 drivers
S_0x5c7c32e190e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e18ec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116cd0 .functor NAND 1, L_0x5c7c33116c20, L_0x5c7c33116c20, C4<1>, C4<1>;
v0x5c7c32e19350_0 .net "in_a", 0 0, L_0x5c7c33116c20;  alias, 1 drivers
v0x5c7c32e19410_0 .net "in_b", 0 0, L_0x5c7c33116c20;  alias, 1 drivers
v0x5c7c32e19560_0 .net "out", 0 0, L_0x5c7c33116cd0;  alias, 1 drivers
S_0x5c7c32e1a8e0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32e02730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e202d0_0 .net "branch1_out", 0 0, L_0x5c7c33116f60;  1 drivers
v0x5c7c32e20400_0 .net "branch2_out", 0 0, L_0x5c7c331171f0;  1 drivers
v0x5c7c32e20550_0 .net "in_a", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e20730_0 .net "in_b", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e208e0_0 .net "out", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e20980_0 .net "temp1_out", 0 0, L_0x5c7c33116eb0;  1 drivers
v0x5c7c32e20a20_0 .net "temp2_out", 0 0, L_0x5c7c33117140;  1 drivers
v0x5c7c32e20ac0_0 .net "temp3_out", 0 0, L_0x5c7c331173d0;  1 drivers
S_0x5c7c32e1aa70 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e1a8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e1bb10_0 .net "in_a", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e1bbb0_0 .net "in_b", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e1bc70_0 .net "out", 0 0, L_0x5c7c33116eb0;  alias, 1 drivers
v0x5c7c32e1bd90_0 .net "temp_out", 0 0, L_0x5c7c32e194f0;  1 drivers
S_0x5c7c32e1ac90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e1aa70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e194f0 .functor NAND 1, L_0x5c7c33115250, L_0x5c7c33115250, C4<1>, C4<1>;
v0x5c7c32e1af00_0 .net "in_a", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e1b050_0 .net "in_b", 0 0, L_0x5c7c33115250;  alias, 1 drivers
v0x5c7c32e1b110_0 .net "out", 0 0, L_0x5c7c32e194f0;  alias, 1 drivers
S_0x5c7c32e1b240 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e1aa70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e1b960_0 .net "in_a", 0 0, L_0x5c7c32e194f0;  alias, 1 drivers
v0x5c7c32e1ba00_0 .net "out", 0 0, L_0x5c7c33116eb0;  alias, 1 drivers
S_0x5c7c32e1b410 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e1b240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116eb0 .functor NAND 1, L_0x5c7c32e194f0, L_0x5c7c32e194f0, C4<1>, C4<1>;
v0x5c7c32e1b680_0 .net "in_a", 0 0, L_0x5c7c32e194f0;  alias, 1 drivers
v0x5c7c32e1b770_0 .net "in_b", 0 0, L_0x5c7c32e194f0;  alias, 1 drivers
v0x5c7c32e1b860_0 .net "out", 0 0, L_0x5c7c33116eb0;  alias, 1 drivers
S_0x5c7c32e1bf00 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e1a8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e1cf30_0 .net "in_a", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e1cfd0_0 .net "in_b", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e1d090_0 .net "out", 0 0, L_0x5c7c33117140;  alias, 1 drivers
v0x5c7c32e1d1b0_0 .net "temp_out", 0 0, L_0x5c7c32e1ed50;  1 drivers
S_0x5c7c32e1c0e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e1bf00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e1ed50 .functor NAND 1, L_0x5c7c331163a0, L_0x5c7c331163a0, C4<1>, C4<1>;
v0x5c7c32e1c350_0 .net "in_a", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e1c4a0_0 .net "in_b", 0 0, L_0x5c7c331163a0;  alias, 1 drivers
v0x5c7c32e1c560_0 .net "out", 0 0, L_0x5c7c32e1ed50;  alias, 1 drivers
S_0x5c7c32e1c660 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e1bf00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e1cd80_0 .net "in_a", 0 0, L_0x5c7c32e1ed50;  alias, 1 drivers
v0x5c7c32e1ce20_0 .net "out", 0 0, L_0x5c7c33117140;  alias, 1 drivers
S_0x5c7c32e1c830 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e1c660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117140 .functor NAND 1, L_0x5c7c32e1ed50, L_0x5c7c32e1ed50, C4<1>, C4<1>;
v0x5c7c32e1caa0_0 .net "in_a", 0 0, L_0x5c7c32e1ed50;  alias, 1 drivers
v0x5c7c32e1cb90_0 .net "in_b", 0 0, L_0x5c7c32e1ed50;  alias, 1 drivers
v0x5c7c32e1cc80_0 .net "out", 0 0, L_0x5c7c33117140;  alias, 1 drivers
S_0x5c7c32e1d320 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e1a8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e1e360_0 .net "in_a", 0 0, L_0x5c7c33116f60;  alias, 1 drivers
v0x5c7c32e1e430_0 .net "in_b", 0 0, L_0x5c7c331171f0;  alias, 1 drivers
v0x5c7c32e1e500_0 .net "out", 0 0, L_0x5c7c331173d0;  alias, 1 drivers
v0x5c7c32e1e620_0 .net "temp_out", 0 0, L_0x5c7c32e1f6c0;  1 drivers
S_0x5c7c32e1d500 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e1d320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e1f6c0 .functor NAND 1, L_0x5c7c33116f60, L_0x5c7c331171f0, C4<1>, C4<1>;
v0x5c7c32e1d750_0 .net "in_a", 0 0, L_0x5c7c33116f60;  alias, 1 drivers
v0x5c7c32e1d830_0 .net "in_b", 0 0, L_0x5c7c331171f0;  alias, 1 drivers
v0x5c7c32e1d8f0_0 .net "out", 0 0, L_0x5c7c32e1f6c0;  alias, 1 drivers
S_0x5c7c32e1da40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e1d320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e1e1b0_0 .net "in_a", 0 0, L_0x5c7c32e1f6c0;  alias, 1 drivers
v0x5c7c32e1e250_0 .net "out", 0 0, L_0x5c7c331173d0;  alias, 1 drivers
S_0x5c7c32e1dc60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e1da40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331173d0 .functor NAND 1, L_0x5c7c32e1f6c0, L_0x5c7c32e1f6c0, C4<1>, C4<1>;
v0x5c7c32e1ded0_0 .net "in_a", 0 0, L_0x5c7c32e1f6c0;  alias, 1 drivers
v0x5c7c32e1dfc0_0 .net "in_b", 0 0, L_0x5c7c32e1f6c0;  alias, 1 drivers
v0x5c7c32e1e0b0_0 .net "out", 0 0, L_0x5c7c331173d0;  alias, 1 drivers
S_0x5c7c32e1e770 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e1a8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e1eea0_0 .net "in_a", 0 0, L_0x5c7c33116eb0;  alias, 1 drivers
v0x5c7c32e1ef40_0 .net "out", 0 0, L_0x5c7c33116f60;  alias, 1 drivers
S_0x5c7c32e1e940 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e1e770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33116f60 .functor NAND 1, L_0x5c7c33116eb0, L_0x5c7c33116eb0, C4<1>, C4<1>;
v0x5c7c32e1ebb0_0 .net "in_a", 0 0, L_0x5c7c33116eb0;  alias, 1 drivers
v0x5c7c32e1ec70_0 .net "in_b", 0 0, L_0x5c7c33116eb0;  alias, 1 drivers
v0x5c7c32e1edc0_0 .net "out", 0 0, L_0x5c7c33116f60;  alias, 1 drivers
S_0x5c7c32e1f040 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e1a8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e1f810_0 .net "in_a", 0 0, L_0x5c7c33117140;  alias, 1 drivers
v0x5c7c32e1f8b0_0 .net "out", 0 0, L_0x5c7c331171f0;  alias, 1 drivers
S_0x5c7c32e1f2b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e1f040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331171f0 .functor NAND 1, L_0x5c7c33117140, L_0x5c7c33117140, C4<1>, C4<1>;
v0x5c7c32e1f520_0 .net "in_a", 0 0, L_0x5c7c33117140;  alias, 1 drivers
v0x5c7c32e1f5e0_0 .net "in_b", 0 0, L_0x5c7c33117140;  alias, 1 drivers
v0x5c7c32e1f730_0 .net "out", 0 0, L_0x5c7c331171f0;  alias, 1 drivers
S_0x5c7c32e1f9b0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e1a8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e20150_0 .net "in_a", 0 0, L_0x5c7c331173d0;  alias, 1 drivers
v0x5c7c32e201f0_0 .net "out", 0 0, L_0x5c7c33117480;  alias, 1 drivers
S_0x5c7c32e1fbd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e1f9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117480 .functor NAND 1, L_0x5c7c331173d0, L_0x5c7c331173d0, C4<1>, C4<1>;
v0x5c7c32e1fe40_0 .net "in_a", 0 0, L_0x5c7c331173d0;  alias, 1 drivers
v0x5c7c32e1ff00_0 .net "in_b", 0 0, L_0x5c7c331173d0;  alias, 1 drivers
v0x5c7c32e20050_0 .net "out", 0 0, L_0x5c7c33117480;  alias, 1 drivers
S_0x5c7c32e21120 .scope module, "fa_gate4" "FullAdder" 2 9, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32e3f550_0 .net "a", 0 0, L_0x5c7c33119bc0;  1 drivers
v0x5c7c32e3f5f0_0 .net "b", 0 0, L_0x5c7c33119c60;  1 drivers
v0x5c7c32e3f6b0_0 .net "c", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e3f750_0 .net "carry", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e3f7f0_0 .net "sum", 0 0, L_0x5c7c33119270;  1 drivers
v0x5c7c32e3f890_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c331177f0;  1 drivers
v0x5c7c32e3f930_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33118940;  1 drivers
v0x5c7c32e3f9d0_0 .net "tmp_sum_out", 0 0, L_0x5c7c33118340;  1 drivers
S_0x5c7c32e21380 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32e21120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e2cf00_0 .net "a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e2d0b0_0 .net "b", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e2d280_0 .net "carry", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e2d320_0 .net "sum", 0 0, L_0x5c7c33118340;  alias, 1 drivers
S_0x5c7c32e215f0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e21380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e226e0_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e227b0_0 .net "in_b", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e22880_0 .net "out", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e229a0_0 .net "temp_out", 0 0, L_0x5c7c33117760;  1 drivers
S_0x5c7c32e21860 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e215f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117760 .functor NAND 1, L_0x5c7c33119bc0, L_0x5c7c33119c60, C4<1>, C4<1>;
v0x5c7c32e21ad0_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e21bb0_0 .net "in_b", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e21c70_0 .net "out", 0 0, L_0x5c7c33117760;  alias, 1 drivers
S_0x5c7c32e21dc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e215f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e22530_0 .net "in_a", 0 0, L_0x5c7c33117760;  alias, 1 drivers
v0x5c7c32e225d0_0 .net "out", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
S_0x5c7c32e21fe0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e21dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331177f0 .functor NAND 1, L_0x5c7c33117760, L_0x5c7c33117760, C4<1>, C4<1>;
v0x5c7c32e22250_0 .net "in_a", 0 0, L_0x5c7c33117760;  alias, 1 drivers
v0x5c7c32e22340_0 .net "in_b", 0 0, L_0x5c7c33117760;  alias, 1 drivers
v0x5c7c32e22430_0 .net "out", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
S_0x5c7c32e22a60 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e21380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e2c820_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e2c8c0_0 .net "in_b", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e2c980_0 .net "out", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e2ca20_0 .net "temp_a_and_out", 0 0, L_0x5c7c33117a00;  1 drivers
v0x5c7c32e2cbd0_0 .net "temp_a_out", 0 0, L_0x5c7c331178a0;  1 drivers
v0x5c7c32e2cc70_0 .net "temp_b_and_out", 0 0, L_0x5c7c33117c10;  1 drivers
v0x5c7c32e2ce20_0 .net "temp_b_out", 0 0, L_0x5c7c33117ab0;  1 drivers
S_0x5c7c32e22c40 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e22a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e23d00_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e23da0_0 .net "in_b", 0 0, L_0x5c7c331178a0;  alias, 1 drivers
v0x5c7c32e23e90_0 .net "out", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
v0x5c7c32e23fb0_0 .net "temp_out", 0 0, L_0x5c7c33117950;  1 drivers
S_0x5c7c32e22eb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e22c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117950 .functor NAND 1, L_0x5c7c33119bc0, L_0x5c7c331178a0, C4<1>, C4<1>;
v0x5c7c32e23120_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e23230_0 .net "in_b", 0 0, L_0x5c7c331178a0;  alias, 1 drivers
v0x5c7c32e232f0_0 .net "out", 0 0, L_0x5c7c33117950;  alias, 1 drivers
S_0x5c7c32e23410 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e22c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e23b50_0 .net "in_a", 0 0, L_0x5c7c33117950;  alias, 1 drivers
v0x5c7c32e23bf0_0 .net "out", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
S_0x5c7c32e23630 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e23410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117a00 .functor NAND 1, L_0x5c7c33117950, L_0x5c7c33117950, C4<1>, C4<1>;
v0x5c7c32e238a0_0 .net "in_a", 0 0, L_0x5c7c33117950;  alias, 1 drivers
v0x5c7c32e23960_0 .net "in_b", 0 0, L_0x5c7c33117950;  alias, 1 drivers
v0x5c7c32e23a50_0 .net "out", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
S_0x5c7c32e24070 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e22a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e250a0_0 .net "in_a", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e25140_0 .net "in_b", 0 0, L_0x5c7c33117ab0;  alias, 1 drivers
v0x5c7c32e25230_0 .net "out", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
v0x5c7c32e25350_0 .net "temp_out", 0 0, L_0x5c7c33117b60;  1 drivers
S_0x5c7c32e24250 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e24070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117b60 .functor NAND 1, L_0x5c7c33119c60, L_0x5c7c33117ab0, C4<1>, C4<1>;
v0x5c7c32e244c0_0 .net "in_a", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e245d0_0 .net "in_b", 0 0, L_0x5c7c33117ab0;  alias, 1 drivers
v0x5c7c32e24690_0 .net "out", 0 0, L_0x5c7c33117b60;  alias, 1 drivers
S_0x5c7c32e247b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e24070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e24ef0_0 .net "in_a", 0 0, L_0x5c7c33117b60;  alias, 1 drivers
v0x5c7c32e24f90_0 .net "out", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
S_0x5c7c32e249d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e247b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117c10 .functor NAND 1, L_0x5c7c33117b60, L_0x5c7c33117b60, C4<1>, C4<1>;
v0x5c7c32e24c40_0 .net "in_a", 0 0, L_0x5c7c33117b60;  alias, 1 drivers
v0x5c7c32e24d00_0 .net "in_b", 0 0, L_0x5c7c33117b60;  alias, 1 drivers
v0x5c7c32e24df0_0 .net "out", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
S_0x5c7c32e254a0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e22a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e25be0_0 .net "in_a", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e25c80_0 .net "out", 0 0, L_0x5c7c331178a0;  alias, 1 drivers
S_0x5c7c32e25670 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e254a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331178a0 .functor NAND 1, L_0x5c7c33119c60, L_0x5c7c33119c60, C4<1>, C4<1>;
v0x5c7c32e258c0_0 .net "in_a", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e25a10_0 .net "in_b", 0 0, L_0x5c7c33119c60;  alias, 1 drivers
v0x5c7c32e25ad0_0 .net "out", 0 0, L_0x5c7c331178a0;  alias, 1 drivers
S_0x5c7c32e25d80 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e22a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e26500_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e265a0_0 .net "out", 0 0, L_0x5c7c33117ab0;  alias, 1 drivers
S_0x5c7c32e25fa0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e25d80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117ab0 .functor NAND 1, L_0x5c7c33119bc0, L_0x5c7c33119bc0, C4<1>, C4<1>;
v0x5c7c32e26210_0 .net "in_a", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e26360_0 .net "in_b", 0 0, L_0x5c7c33119bc0;  alias, 1 drivers
v0x5c7c32e26420_0 .net "out", 0 0, L_0x5c7c33117ab0;  alias, 1 drivers
S_0x5c7c32e266a0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e22a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e2c170_0 .net "branch1_out", 0 0, L_0x5c7c33117e20;  1 drivers
v0x5c7c32e2c2a0_0 .net "branch2_out", 0 0, L_0x5c7c331180b0;  1 drivers
v0x5c7c32e2c3f0_0 .net "in_a", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
v0x5c7c32e2c4c0_0 .net "in_b", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
v0x5c7c32e2c560_0 .net "out", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e2c600_0 .net "temp1_out", 0 0, L_0x5c7c33117d70;  1 drivers
v0x5c7c32e2c6a0_0 .net "temp2_out", 0 0, L_0x5c7c33118000;  1 drivers
v0x5c7c32e2c740_0 .net "temp3_out", 0 0, L_0x5c7c33118290;  1 drivers
S_0x5c7c32e26920 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e266a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e279b0_0 .net "in_a", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
v0x5c7c32e27a50_0 .net "in_b", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
v0x5c7c32e27b10_0 .net "out", 0 0, L_0x5c7c33117d70;  alias, 1 drivers
v0x5c7c32e27c30_0 .net "temp_out", 0 0, L_0x5c7c33117cc0;  1 drivers
S_0x5c7c32e26b90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e26920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117cc0 .functor NAND 1, L_0x5c7c33117a00, L_0x5c7c33117a00, C4<1>, C4<1>;
v0x5c7c32e26e00_0 .net "in_a", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
v0x5c7c32e26ec0_0 .net "in_b", 0 0, L_0x5c7c33117a00;  alias, 1 drivers
v0x5c7c32e27010_0 .net "out", 0 0, L_0x5c7c33117cc0;  alias, 1 drivers
S_0x5c7c32e27110 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e26920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e27800_0 .net "in_a", 0 0, L_0x5c7c33117cc0;  alias, 1 drivers
v0x5c7c32e278a0_0 .net "out", 0 0, L_0x5c7c33117d70;  alias, 1 drivers
S_0x5c7c32e272e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e27110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117d70 .functor NAND 1, L_0x5c7c33117cc0, L_0x5c7c33117cc0, C4<1>, C4<1>;
v0x5c7c32e27550_0 .net "in_a", 0 0, L_0x5c7c33117cc0;  alias, 1 drivers
v0x5c7c32e27610_0 .net "in_b", 0 0, L_0x5c7c33117cc0;  alias, 1 drivers
v0x5c7c32e27700_0 .net "out", 0 0, L_0x5c7c33117d70;  alias, 1 drivers
S_0x5c7c32e27da0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e266a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e28dd0_0 .net "in_a", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
v0x5c7c32e28e70_0 .net "in_b", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
v0x5c7c32e28f30_0 .net "out", 0 0, L_0x5c7c33118000;  alias, 1 drivers
v0x5c7c32e29050_0 .net "temp_out", 0 0, L_0x5c7c32e2abf0;  1 drivers
S_0x5c7c32e27f80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e27da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e2abf0 .functor NAND 1, L_0x5c7c33117c10, L_0x5c7c33117c10, C4<1>, C4<1>;
v0x5c7c32e281f0_0 .net "in_a", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
v0x5c7c32e282b0_0 .net "in_b", 0 0, L_0x5c7c33117c10;  alias, 1 drivers
v0x5c7c32e28400_0 .net "out", 0 0, L_0x5c7c32e2abf0;  alias, 1 drivers
S_0x5c7c32e28500 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e27da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e28c20_0 .net "in_a", 0 0, L_0x5c7c32e2abf0;  alias, 1 drivers
v0x5c7c32e28cc0_0 .net "out", 0 0, L_0x5c7c33118000;  alias, 1 drivers
S_0x5c7c32e286d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e28500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118000 .functor NAND 1, L_0x5c7c32e2abf0, L_0x5c7c32e2abf0, C4<1>, C4<1>;
v0x5c7c32e28940_0 .net "in_a", 0 0, L_0x5c7c32e2abf0;  alias, 1 drivers
v0x5c7c32e28a30_0 .net "in_b", 0 0, L_0x5c7c32e2abf0;  alias, 1 drivers
v0x5c7c32e28b20_0 .net "out", 0 0, L_0x5c7c33118000;  alias, 1 drivers
S_0x5c7c32e291c0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e266a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e2a200_0 .net "in_a", 0 0, L_0x5c7c33117e20;  alias, 1 drivers
v0x5c7c32e2a2d0_0 .net "in_b", 0 0, L_0x5c7c331180b0;  alias, 1 drivers
v0x5c7c32e2a3a0_0 .net "out", 0 0, L_0x5c7c33118290;  alias, 1 drivers
v0x5c7c32e2a4c0_0 .net "temp_out", 0 0, L_0x5c7c32e2b560;  1 drivers
S_0x5c7c32e293a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e291c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e2b560 .functor NAND 1, L_0x5c7c33117e20, L_0x5c7c331180b0, C4<1>, C4<1>;
v0x5c7c32e295f0_0 .net "in_a", 0 0, L_0x5c7c33117e20;  alias, 1 drivers
v0x5c7c32e296d0_0 .net "in_b", 0 0, L_0x5c7c331180b0;  alias, 1 drivers
v0x5c7c32e29790_0 .net "out", 0 0, L_0x5c7c32e2b560;  alias, 1 drivers
S_0x5c7c32e298e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e291c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e2a050_0 .net "in_a", 0 0, L_0x5c7c32e2b560;  alias, 1 drivers
v0x5c7c32e2a0f0_0 .net "out", 0 0, L_0x5c7c33118290;  alias, 1 drivers
S_0x5c7c32e29b00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e298e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118290 .functor NAND 1, L_0x5c7c32e2b560, L_0x5c7c32e2b560, C4<1>, C4<1>;
v0x5c7c32e29d70_0 .net "in_a", 0 0, L_0x5c7c32e2b560;  alias, 1 drivers
v0x5c7c32e29e60_0 .net "in_b", 0 0, L_0x5c7c32e2b560;  alias, 1 drivers
v0x5c7c32e29f50_0 .net "out", 0 0, L_0x5c7c33118290;  alias, 1 drivers
S_0x5c7c32e2a610 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e266a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e2ad40_0 .net "in_a", 0 0, L_0x5c7c33117d70;  alias, 1 drivers
v0x5c7c32e2ade0_0 .net "out", 0 0, L_0x5c7c33117e20;  alias, 1 drivers
S_0x5c7c32e2a7e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e2a610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33117e20 .functor NAND 1, L_0x5c7c33117d70, L_0x5c7c33117d70, C4<1>, C4<1>;
v0x5c7c32e2aa50_0 .net "in_a", 0 0, L_0x5c7c33117d70;  alias, 1 drivers
v0x5c7c32e2ab10_0 .net "in_b", 0 0, L_0x5c7c33117d70;  alias, 1 drivers
v0x5c7c32e2ac60_0 .net "out", 0 0, L_0x5c7c33117e20;  alias, 1 drivers
S_0x5c7c32e2aee0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e266a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e2b6b0_0 .net "in_a", 0 0, L_0x5c7c33118000;  alias, 1 drivers
v0x5c7c32e2b750_0 .net "out", 0 0, L_0x5c7c331180b0;  alias, 1 drivers
S_0x5c7c32e2b150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e2aee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331180b0 .functor NAND 1, L_0x5c7c33118000, L_0x5c7c33118000, C4<1>, C4<1>;
v0x5c7c32e2b3c0_0 .net "in_a", 0 0, L_0x5c7c33118000;  alias, 1 drivers
v0x5c7c32e2b480_0 .net "in_b", 0 0, L_0x5c7c33118000;  alias, 1 drivers
v0x5c7c32e2b5d0_0 .net "out", 0 0, L_0x5c7c331180b0;  alias, 1 drivers
S_0x5c7c32e2b850 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e266a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e2bff0_0 .net "in_a", 0 0, L_0x5c7c33118290;  alias, 1 drivers
v0x5c7c32e2c090_0 .net "out", 0 0, L_0x5c7c33118340;  alias, 1 drivers
S_0x5c7c32e2ba70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e2b850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118340 .functor NAND 1, L_0x5c7c33118290, L_0x5c7c33118290, C4<1>, C4<1>;
v0x5c7c32e2bce0_0 .net "in_a", 0 0, L_0x5c7c33118290;  alias, 1 drivers
v0x5c7c32e2bda0_0 .net "in_b", 0 0, L_0x5c7c33118290;  alias, 1 drivers
v0x5c7c32e2bef0_0 .net "out", 0 0, L_0x5c7c33118340;  alias, 1 drivers
S_0x5c7c32e2d400 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32e21120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e38f20_0 .net "a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e38fc0_0 .net "b", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e39080_0 .net "carry", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e39120_0 .net "sum", 0 0, L_0x5c7c33119270;  alias, 1 drivers
S_0x5c7c32e2d620 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e2d400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e2e5c0_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e2e660_0 .net "in_b", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e2e720_0 .net "out", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e2e840_0 .net "temp_out", 0 0, L_0x5c7c32e2be80;  1 drivers
S_0x5c7c32e2d7d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e2d620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e2be80 .functor NAND 1, L_0x5c7c33118340, L_0x5c7c33117480, C4<1>, C4<1>;
v0x5c7c32e2da40_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e2db00_0 .net "in_b", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e2dbc0_0 .net "out", 0 0, L_0x5c7c32e2be80;  alias, 1 drivers
S_0x5c7c32e2dcf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e2d620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e2e410_0 .net "in_a", 0 0, L_0x5c7c32e2be80;  alias, 1 drivers
v0x5c7c32e2e4b0_0 .net "out", 0 0, L_0x5c7c33118940;  alias, 1 drivers
S_0x5c7c32e2dec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e2dcf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118940 .functor NAND 1, L_0x5c7c32e2be80, L_0x5c7c32e2be80, C4<1>, C4<1>;
v0x5c7c32e2e130_0 .net "in_a", 0 0, L_0x5c7c32e2be80;  alias, 1 drivers
v0x5c7c32e2e220_0 .net "in_b", 0 0, L_0x5c7c32e2be80;  alias, 1 drivers
v0x5c7c32e2e310_0 .net "out", 0 0, L_0x5c7c33118940;  alias, 1 drivers
S_0x5c7c32e2e9b0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e2d400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e38840_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e388e0_0 .net "in_b", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e389a0_0 .net "out", 0 0, L_0x5c7c33119270;  alias, 1 drivers
v0x5c7c32e38a40_0 .net "temp_a_and_out", 0 0, L_0x5c7c33118b50;  1 drivers
v0x5c7c32e38bf0_0 .net "temp_a_out", 0 0, L_0x5c7c331189f0;  1 drivers
v0x5c7c32e38c90_0 .net "temp_b_and_out", 0 0, L_0x5c7c33118d60;  1 drivers
v0x5c7c32e38e40_0 .net "temp_b_out", 0 0, L_0x5c7c33118c00;  1 drivers
S_0x5c7c32e2eb90 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e2e9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e2fc30_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e2fde0_0 .net "in_b", 0 0, L_0x5c7c331189f0;  alias, 1 drivers
v0x5c7c32e2fed0_0 .net "out", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
v0x5c7c32e2fff0_0 .net "temp_out", 0 0, L_0x5c7c33118aa0;  1 drivers
S_0x5c7c32e2ee00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e2eb90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118aa0 .functor NAND 1, L_0x5c7c33118340, L_0x5c7c331189f0, C4<1>, C4<1>;
v0x5c7c32e2f070_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e2f130_0 .net "in_b", 0 0, L_0x5c7c331189f0;  alias, 1 drivers
v0x5c7c32e2f1f0_0 .net "out", 0 0, L_0x5c7c33118aa0;  alias, 1 drivers
S_0x5c7c32e2f310 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e2eb90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e2fa80_0 .net "in_a", 0 0, L_0x5c7c33118aa0;  alias, 1 drivers
v0x5c7c32e2fb20_0 .net "out", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
S_0x5c7c32e2f530 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e2f310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118b50 .functor NAND 1, L_0x5c7c33118aa0, L_0x5c7c33118aa0, C4<1>, C4<1>;
v0x5c7c32e2f7a0_0 .net "in_a", 0 0, L_0x5c7c33118aa0;  alias, 1 drivers
v0x5c7c32e2f890_0 .net "in_b", 0 0, L_0x5c7c33118aa0;  alias, 1 drivers
v0x5c7c32e2f980_0 .net "out", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
S_0x5c7c32e300b0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e2e9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e310c0_0 .net "in_a", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e31160_0 .net "in_b", 0 0, L_0x5c7c33118c00;  alias, 1 drivers
v0x5c7c32e31250_0 .net "out", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
v0x5c7c32e31370_0 .net "temp_out", 0 0, L_0x5c7c33118cb0;  1 drivers
S_0x5c7c32e30290 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e300b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118cb0 .functor NAND 1, L_0x5c7c33117480, L_0x5c7c33118c00, C4<1>, C4<1>;
v0x5c7c32e30500_0 .net "in_a", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e305c0_0 .net "in_b", 0 0, L_0x5c7c33118c00;  alias, 1 drivers
v0x5c7c32e30680_0 .net "out", 0 0, L_0x5c7c33118cb0;  alias, 1 drivers
S_0x5c7c32e307a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e300b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e30f10_0 .net "in_a", 0 0, L_0x5c7c33118cb0;  alias, 1 drivers
v0x5c7c32e30fb0_0 .net "out", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
S_0x5c7c32e309c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e307a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118d60 .functor NAND 1, L_0x5c7c33118cb0, L_0x5c7c33118cb0, C4<1>, C4<1>;
v0x5c7c32e30c30_0 .net "in_a", 0 0, L_0x5c7c33118cb0;  alias, 1 drivers
v0x5c7c32e30d20_0 .net "in_b", 0 0, L_0x5c7c33118cb0;  alias, 1 drivers
v0x5c7c32e30e10_0 .net "out", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
S_0x5c7c32e314c0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e2e9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e31cd0_0 .net "in_a", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e31d70_0 .net "out", 0 0, L_0x5c7c331189f0;  alias, 1 drivers
S_0x5c7c32e31690 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e314c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331189f0 .functor NAND 1, L_0x5c7c33117480, L_0x5c7c33117480, C4<1>, C4<1>;
v0x5c7c32e318e0_0 .net "in_a", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e31ab0_0 .net "in_b", 0 0, L_0x5c7c33117480;  alias, 1 drivers
v0x5c7c32e31b70_0 .net "out", 0 0, L_0x5c7c331189f0;  alias, 1 drivers
S_0x5c7c32e31e70 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e2e9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e325b0_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e32650_0 .net "out", 0 0, L_0x5c7c33118c00;  alias, 1 drivers
S_0x5c7c32e32090 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e31e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118c00 .functor NAND 1, L_0x5c7c33118340, L_0x5c7c33118340, C4<1>, C4<1>;
v0x5c7c32e32300_0 .net "in_a", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e323c0_0 .net "in_b", 0 0, L_0x5c7c33118340;  alias, 1 drivers
v0x5c7c32e32480_0 .net "out", 0 0, L_0x5c7c33118c00;  alias, 1 drivers
S_0x5c7c32e32750 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e2e9b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e38190_0 .net "branch1_out", 0 0, L_0x5c7c33118f70;  1 drivers
v0x5c7c32e382c0_0 .net "branch2_out", 0 0, L_0x5c7c331190f0;  1 drivers
v0x5c7c32e38410_0 .net "in_a", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
v0x5c7c32e384e0_0 .net "in_b", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
v0x5c7c32e38580_0 .net "out", 0 0, L_0x5c7c33119270;  alias, 1 drivers
v0x5c7c32e38620_0 .net "temp1_out", 0 0, L_0x5c7c33118ec0;  1 drivers
v0x5c7c32e386c0_0 .net "temp2_out", 0 0, L_0x5c7c33119040;  1 drivers
v0x5c7c32e38760_0 .net "temp3_out", 0 0, L_0x5c7c331191c0;  1 drivers
S_0x5c7c32e329d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e32750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e339d0_0 .net "in_a", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
v0x5c7c32e33a70_0 .net "in_b", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
v0x5c7c32e33b30_0 .net "out", 0 0, L_0x5c7c33118ec0;  alias, 1 drivers
v0x5c7c32e33c50_0 .net "temp_out", 0 0, L_0x5c7c33118e10;  1 drivers
S_0x5c7c32e32c40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e329d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118e10 .functor NAND 1, L_0x5c7c33118b50, L_0x5c7c33118b50, C4<1>, C4<1>;
v0x5c7c32e32eb0_0 .net "in_a", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
v0x5c7c32e32f70_0 .net "in_b", 0 0, L_0x5c7c33118b50;  alias, 1 drivers
v0x5c7c32e33030_0 .net "out", 0 0, L_0x5c7c33118e10;  alias, 1 drivers
S_0x5c7c32e33130 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e329d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e33820_0 .net "in_a", 0 0, L_0x5c7c33118e10;  alias, 1 drivers
v0x5c7c32e338c0_0 .net "out", 0 0, L_0x5c7c33118ec0;  alias, 1 drivers
S_0x5c7c32e33300 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e33130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118ec0 .functor NAND 1, L_0x5c7c33118e10, L_0x5c7c33118e10, C4<1>, C4<1>;
v0x5c7c32e33570_0 .net "in_a", 0 0, L_0x5c7c33118e10;  alias, 1 drivers
v0x5c7c32e33630_0 .net "in_b", 0 0, L_0x5c7c33118e10;  alias, 1 drivers
v0x5c7c32e33720_0 .net "out", 0 0, L_0x5c7c33118ec0;  alias, 1 drivers
S_0x5c7c32e33dc0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e32750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e34df0_0 .net "in_a", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
v0x5c7c32e34e90_0 .net "in_b", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
v0x5c7c32e34f50_0 .net "out", 0 0, L_0x5c7c33119040;  alias, 1 drivers
v0x5c7c32e35070_0 .net "temp_out", 0 0, L_0x5c7c32e36c10;  1 drivers
S_0x5c7c32e33fa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e33dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e36c10 .functor NAND 1, L_0x5c7c33118d60, L_0x5c7c33118d60, C4<1>, C4<1>;
v0x5c7c32e34210_0 .net "in_a", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
v0x5c7c32e342d0_0 .net "in_b", 0 0, L_0x5c7c33118d60;  alias, 1 drivers
v0x5c7c32e34420_0 .net "out", 0 0, L_0x5c7c32e36c10;  alias, 1 drivers
S_0x5c7c32e34520 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e33dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e34c40_0 .net "in_a", 0 0, L_0x5c7c32e36c10;  alias, 1 drivers
v0x5c7c32e34ce0_0 .net "out", 0 0, L_0x5c7c33119040;  alias, 1 drivers
S_0x5c7c32e346f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e34520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119040 .functor NAND 1, L_0x5c7c32e36c10, L_0x5c7c32e36c10, C4<1>, C4<1>;
v0x5c7c32e34960_0 .net "in_a", 0 0, L_0x5c7c32e36c10;  alias, 1 drivers
v0x5c7c32e34a50_0 .net "in_b", 0 0, L_0x5c7c32e36c10;  alias, 1 drivers
v0x5c7c32e34b40_0 .net "out", 0 0, L_0x5c7c33119040;  alias, 1 drivers
S_0x5c7c32e351e0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e32750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e36220_0 .net "in_a", 0 0, L_0x5c7c33118f70;  alias, 1 drivers
v0x5c7c32e362f0_0 .net "in_b", 0 0, L_0x5c7c331190f0;  alias, 1 drivers
v0x5c7c32e363c0_0 .net "out", 0 0, L_0x5c7c331191c0;  alias, 1 drivers
v0x5c7c32e364e0_0 .net "temp_out", 0 0, L_0x5c7c32e37580;  1 drivers
S_0x5c7c32e353c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e351e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e37580 .functor NAND 1, L_0x5c7c33118f70, L_0x5c7c331190f0, C4<1>, C4<1>;
v0x5c7c32e35610_0 .net "in_a", 0 0, L_0x5c7c33118f70;  alias, 1 drivers
v0x5c7c32e356f0_0 .net "in_b", 0 0, L_0x5c7c331190f0;  alias, 1 drivers
v0x5c7c32e357b0_0 .net "out", 0 0, L_0x5c7c32e37580;  alias, 1 drivers
S_0x5c7c32e35900 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e351e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e36070_0 .net "in_a", 0 0, L_0x5c7c32e37580;  alias, 1 drivers
v0x5c7c32e36110_0 .net "out", 0 0, L_0x5c7c331191c0;  alias, 1 drivers
S_0x5c7c32e35b20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e35900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331191c0 .functor NAND 1, L_0x5c7c32e37580, L_0x5c7c32e37580, C4<1>, C4<1>;
v0x5c7c32e35d90_0 .net "in_a", 0 0, L_0x5c7c32e37580;  alias, 1 drivers
v0x5c7c32e35e80_0 .net "in_b", 0 0, L_0x5c7c32e37580;  alias, 1 drivers
v0x5c7c32e35f70_0 .net "out", 0 0, L_0x5c7c331191c0;  alias, 1 drivers
S_0x5c7c32e36630 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e32750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e36d60_0 .net "in_a", 0 0, L_0x5c7c33118ec0;  alias, 1 drivers
v0x5c7c32e36e00_0 .net "out", 0 0, L_0x5c7c33118f70;  alias, 1 drivers
S_0x5c7c32e36800 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e36630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33118f70 .functor NAND 1, L_0x5c7c33118ec0, L_0x5c7c33118ec0, C4<1>, C4<1>;
v0x5c7c32e36a70_0 .net "in_a", 0 0, L_0x5c7c33118ec0;  alias, 1 drivers
v0x5c7c32e36b30_0 .net "in_b", 0 0, L_0x5c7c33118ec0;  alias, 1 drivers
v0x5c7c32e36c80_0 .net "out", 0 0, L_0x5c7c33118f70;  alias, 1 drivers
S_0x5c7c32e36f00 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e32750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e376d0_0 .net "in_a", 0 0, L_0x5c7c33119040;  alias, 1 drivers
v0x5c7c32e37770_0 .net "out", 0 0, L_0x5c7c331190f0;  alias, 1 drivers
S_0x5c7c32e37170 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e36f00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331190f0 .functor NAND 1, L_0x5c7c33119040, L_0x5c7c33119040, C4<1>, C4<1>;
v0x5c7c32e373e0_0 .net "in_a", 0 0, L_0x5c7c33119040;  alias, 1 drivers
v0x5c7c32e374a0_0 .net "in_b", 0 0, L_0x5c7c33119040;  alias, 1 drivers
v0x5c7c32e375f0_0 .net "out", 0 0, L_0x5c7c331190f0;  alias, 1 drivers
S_0x5c7c32e37870 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e32750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e38010_0 .net "in_a", 0 0, L_0x5c7c331191c0;  alias, 1 drivers
v0x5c7c32e380b0_0 .net "out", 0 0, L_0x5c7c33119270;  alias, 1 drivers
S_0x5c7c32e37a90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e37870;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119270 .functor NAND 1, L_0x5c7c331191c0, L_0x5c7c331191c0, C4<1>, C4<1>;
v0x5c7c32e37d00_0 .net "in_a", 0 0, L_0x5c7c331191c0;  alias, 1 drivers
v0x5c7c32e37dc0_0 .net "in_b", 0 0, L_0x5c7c331191c0;  alias, 1 drivers
v0x5c7c32e37f10_0 .net "out", 0 0, L_0x5c7c33119270;  alias, 1 drivers
S_0x5c7c32e39290 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32e21120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e3ec80_0 .net "branch1_out", 0 0, L_0x5c7c33119500;  1 drivers
v0x5c7c32e3edb0_0 .net "branch2_out", 0 0, L_0x5c7c33119790;  1 drivers
v0x5c7c32e3ef00_0 .net "in_a", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e3f0e0_0 .net "in_b", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e3f290_0 .net "out", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e3f330_0 .net "temp1_out", 0 0, L_0x5c7c33119450;  1 drivers
v0x5c7c32e3f3d0_0 .net "temp2_out", 0 0, L_0x5c7c331196e0;  1 drivers
v0x5c7c32e3f470_0 .net "temp3_out", 0 0, L_0x5c7c33119970;  1 drivers
S_0x5c7c32e39420 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e39290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e3a4c0_0 .net "in_a", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e3a560_0 .net "in_b", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e3a620_0 .net "out", 0 0, L_0x5c7c33119450;  alias, 1 drivers
v0x5c7c32e3a740_0 .net "temp_out", 0 0, L_0x5c7c32e37ea0;  1 drivers
S_0x5c7c32e39640 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e39420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e37ea0 .functor NAND 1, L_0x5c7c331177f0, L_0x5c7c331177f0, C4<1>, C4<1>;
v0x5c7c32e398b0_0 .net "in_a", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e39a00_0 .net "in_b", 0 0, L_0x5c7c331177f0;  alias, 1 drivers
v0x5c7c32e39ac0_0 .net "out", 0 0, L_0x5c7c32e37ea0;  alias, 1 drivers
S_0x5c7c32e39bf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e39420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e3a310_0 .net "in_a", 0 0, L_0x5c7c32e37ea0;  alias, 1 drivers
v0x5c7c32e3a3b0_0 .net "out", 0 0, L_0x5c7c33119450;  alias, 1 drivers
S_0x5c7c32e39dc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e39bf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119450 .functor NAND 1, L_0x5c7c32e37ea0, L_0x5c7c32e37ea0, C4<1>, C4<1>;
v0x5c7c32e3a030_0 .net "in_a", 0 0, L_0x5c7c32e37ea0;  alias, 1 drivers
v0x5c7c32e3a120_0 .net "in_b", 0 0, L_0x5c7c32e37ea0;  alias, 1 drivers
v0x5c7c32e3a210_0 .net "out", 0 0, L_0x5c7c33119450;  alias, 1 drivers
S_0x5c7c32e3a8b0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e39290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e3b8e0_0 .net "in_a", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e3b980_0 .net "in_b", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e3ba40_0 .net "out", 0 0, L_0x5c7c331196e0;  alias, 1 drivers
v0x5c7c32e3bb60_0 .net "temp_out", 0 0, L_0x5c7c32e3d700;  1 drivers
S_0x5c7c32e3aa90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e3a8b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e3d700 .functor NAND 1, L_0x5c7c33118940, L_0x5c7c33118940, C4<1>, C4<1>;
v0x5c7c32e3ad00_0 .net "in_a", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e3ae50_0 .net "in_b", 0 0, L_0x5c7c33118940;  alias, 1 drivers
v0x5c7c32e3af10_0 .net "out", 0 0, L_0x5c7c32e3d700;  alias, 1 drivers
S_0x5c7c32e3b010 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e3a8b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e3b730_0 .net "in_a", 0 0, L_0x5c7c32e3d700;  alias, 1 drivers
v0x5c7c32e3b7d0_0 .net "out", 0 0, L_0x5c7c331196e0;  alias, 1 drivers
S_0x5c7c32e3b1e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e3b010;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331196e0 .functor NAND 1, L_0x5c7c32e3d700, L_0x5c7c32e3d700, C4<1>, C4<1>;
v0x5c7c32e3b450_0 .net "in_a", 0 0, L_0x5c7c32e3d700;  alias, 1 drivers
v0x5c7c32e3b540_0 .net "in_b", 0 0, L_0x5c7c32e3d700;  alias, 1 drivers
v0x5c7c32e3b630_0 .net "out", 0 0, L_0x5c7c331196e0;  alias, 1 drivers
S_0x5c7c32e3bcd0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e39290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e3cd10_0 .net "in_a", 0 0, L_0x5c7c33119500;  alias, 1 drivers
v0x5c7c32e3cde0_0 .net "in_b", 0 0, L_0x5c7c33119790;  alias, 1 drivers
v0x5c7c32e3ceb0_0 .net "out", 0 0, L_0x5c7c33119970;  alias, 1 drivers
v0x5c7c32e3cfd0_0 .net "temp_out", 0 0, L_0x5c7c32e3e070;  1 drivers
S_0x5c7c32e3beb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e3bcd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e3e070 .functor NAND 1, L_0x5c7c33119500, L_0x5c7c33119790, C4<1>, C4<1>;
v0x5c7c32e3c100_0 .net "in_a", 0 0, L_0x5c7c33119500;  alias, 1 drivers
v0x5c7c32e3c1e0_0 .net "in_b", 0 0, L_0x5c7c33119790;  alias, 1 drivers
v0x5c7c32e3c2a0_0 .net "out", 0 0, L_0x5c7c32e3e070;  alias, 1 drivers
S_0x5c7c32e3c3f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e3bcd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e3cb60_0 .net "in_a", 0 0, L_0x5c7c32e3e070;  alias, 1 drivers
v0x5c7c32e3cc00_0 .net "out", 0 0, L_0x5c7c33119970;  alias, 1 drivers
S_0x5c7c32e3c610 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e3c3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119970 .functor NAND 1, L_0x5c7c32e3e070, L_0x5c7c32e3e070, C4<1>, C4<1>;
v0x5c7c32e3c880_0 .net "in_a", 0 0, L_0x5c7c32e3e070;  alias, 1 drivers
v0x5c7c32e3c970_0 .net "in_b", 0 0, L_0x5c7c32e3e070;  alias, 1 drivers
v0x5c7c32e3ca60_0 .net "out", 0 0, L_0x5c7c33119970;  alias, 1 drivers
S_0x5c7c32e3d120 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e39290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e3d850_0 .net "in_a", 0 0, L_0x5c7c33119450;  alias, 1 drivers
v0x5c7c32e3d8f0_0 .net "out", 0 0, L_0x5c7c33119500;  alias, 1 drivers
S_0x5c7c32e3d2f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e3d120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119500 .functor NAND 1, L_0x5c7c33119450, L_0x5c7c33119450, C4<1>, C4<1>;
v0x5c7c32e3d560_0 .net "in_a", 0 0, L_0x5c7c33119450;  alias, 1 drivers
v0x5c7c32e3d620_0 .net "in_b", 0 0, L_0x5c7c33119450;  alias, 1 drivers
v0x5c7c32e3d770_0 .net "out", 0 0, L_0x5c7c33119500;  alias, 1 drivers
S_0x5c7c32e3d9f0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e39290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e3e1c0_0 .net "in_a", 0 0, L_0x5c7c331196e0;  alias, 1 drivers
v0x5c7c32e3e260_0 .net "out", 0 0, L_0x5c7c33119790;  alias, 1 drivers
S_0x5c7c32e3dc60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e3d9f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119790 .functor NAND 1, L_0x5c7c331196e0, L_0x5c7c331196e0, C4<1>, C4<1>;
v0x5c7c32e3ded0_0 .net "in_a", 0 0, L_0x5c7c331196e0;  alias, 1 drivers
v0x5c7c32e3df90_0 .net "in_b", 0 0, L_0x5c7c331196e0;  alias, 1 drivers
v0x5c7c32e3e0e0_0 .net "out", 0 0, L_0x5c7c33119790;  alias, 1 drivers
S_0x5c7c32e3e360 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e39290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e3eb00_0 .net "in_a", 0 0, L_0x5c7c33119970;  alias, 1 drivers
v0x5c7c32e3eba0_0 .net "out", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
S_0x5c7c32e3e580 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e3e360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119a20 .functor NAND 1, L_0x5c7c33119970, L_0x5c7c33119970, C4<1>, C4<1>;
v0x5c7c32e3e7f0_0 .net "in_a", 0 0, L_0x5c7c33119970;  alias, 1 drivers
v0x5c7c32e3e8b0_0 .net "in_b", 0 0, L_0x5c7c33119970;  alias, 1 drivers
v0x5c7c32e3ea00_0 .net "out", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
S_0x5c7c32e3fad0 .scope module, "fa_gate5" "FullAdder" 2 10, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32e5df00_0 .net "a", 0 0, L_0x5c7c3311c280;  1 drivers
v0x5c7c32e5dfa0_0 .net "b", 0 0, L_0x5c7c3311c320;  1 drivers
v0x5c7c32e5e060_0 .net "c", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e5e100_0 .net "carry", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e5e1a0_0 .net "sum", 0 0, L_0x5c7c3311b930;  1 drivers
v0x5c7c32e5e240_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33119d90;  1 drivers
v0x5c7c32e5e2e0_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c3311b000;  1 drivers
v0x5c7c32e5e380_0 .net "tmp_sum_out", 0 0, L_0x5c7c3311aa00;  1 drivers
S_0x5c7c32e3fd30 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32e3fad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e4b8b0_0 .net "a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e4ba60_0 .net "b", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e4bc30_0 .net "carry", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e4bcd0_0 .net "sum", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
S_0x5c7c32e3ffa0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e3fd30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e41090_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e41160_0 .net "in_b", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e41230_0 .net "out", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e41350_0 .net "temp_out", 0 0, L_0x5c7c33119d00;  1 drivers
S_0x5c7c32e40210 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e3ffa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119d00 .functor NAND 1, L_0x5c7c3311c280, L_0x5c7c3311c320, C4<1>, C4<1>;
v0x5c7c32e40480_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e40560_0 .net "in_b", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e40620_0 .net "out", 0 0, L_0x5c7c33119d00;  alias, 1 drivers
S_0x5c7c32e40770 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e3ffa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e40ee0_0 .net "in_a", 0 0, L_0x5c7c33119d00;  alias, 1 drivers
v0x5c7c32e40f80_0 .net "out", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
S_0x5c7c32e40990 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e40770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119d90 .functor NAND 1, L_0x5c7c33119d00, L_0x5c7c33119d00, C4<1>, C4<1>;
v0x5c7c32e40c00_0 .net "in_a", 0 0, L_0x5c7c33119d00;  alias, 1 drivers
v0x5c7c32e40cf0_0 .net "in_b", 0 0, L_0x5c7c33119d00;  alias, 1 drivers
v0x5c7c32e40de0_0 .net "out", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
S_0x5c7c32e41410 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e3fd30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e4b1d0_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e4b270_0 .net "in_b", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e4b330_0 .net "out", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e4b3d0_0 .net "temp_a_and_out", 0 0, L_0x5c7c33119fa0;  1 drivers
v0x5c7c32e4b580_0 .net "temp_a_out", 0 0, L_0x5c7c33119e40;  1 drivers
v0x5c7c32e4b620_0 .net "temp_b_and_out", 0 0, L_0x5c7c3311a1b0;  1 drivers
v0x5c7c32e4b7d0_0 .net "temp_b_out", 0 0, L_0x5c7c3311a050;  1 drivers
S_0x5c7c32e415f0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e41410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e426b0_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e42750_0 .net "in_b", 0 0, L_0x5c7c33119e40;  alias, 1 drivers
v0x5c7c32e42840_0 .net "out", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
v0x5c7c32e42960_0 .net "temp_out", 0 0, L_0x5c7c33119ef0;  1 drivers
S_0x5c7c32e41860 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e415f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119ef0 .functor NAND 1, L_0x5c7c3311c280, L_0x5c7c33119e40, C4<1>, C4<1>;
v0x5c7c32e41ad0_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e41be0_0 .net "in_b", 0 0, L_0x5c7c33119e40;  alias, 1 drivers
v0x5c7c32e41ca0_0 .net "out", 0 0, L_0x5c7c33119ef0;  alias, 1 drivers
S_0x5c7c32e41dc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e415f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e42500_0 .net "in_a", 0 0, L_0x5c7c33119ef0;  alias, 1 drivers
v0x5c7c32e425a0_0 .net "out", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
S_0x5c7c32e41fe0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e41dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119fa0 .functor NAND 1, L_0x5c7c33119ef0, L_0x5c7c33119ef0, C4<1>, C4<1>;
v0x5c7c32e42250_0 .net "in_a", 0 0, L_0x5c7c33119ef0;  alias, 1 drivers
v0x5c7c32e42310_0 .net "in_b", 0 0, L_0x5c7c33119ef0;  alias, 1 drivers
v0x5c7c32e42400_0 .net "out", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
S_0x5c7c32e42a20 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e41410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e43a50_0 .net "in_a", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e43af0_0 .net "in_b", 0 0, L_0x5c7c3311a050;  alias, 1 drivers
v0x5c7c32e43be0_0 .net "out", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
v0x5c7c32e43d00_0 .net "temp_out", 0 0, L_0x5c7c3311a100;  1 drivers
S_0x5c7c32e42c00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e42a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a100 .functor NAND 1, L_0x5c7c3311c320, L_0x5c7c3311a050, C4<1>, C4<1>;
v0x5c7c32e42e70_0 .net "in_a", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e42f80_0 .net "in_b", 0 0, L_0x5c7c3311a050;  alias, 1 drivers
v0x5c7c32e43040_0 .net "out", 0 0, L_0x5c7c3311a100;  alias, 1 drivers
S_0x5c7c32e43160 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e42a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e438a0_0 .net "in_a", 0 0, L_0x5c7c3311a100;  alias, 1 drivers
v0x5c7c32e43940_0 .net "out", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
S_0x5c7c32e43380 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e43160;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a1b0 .functor NAND 1, L_0x5c7c3311a100, L_0x5c7c3311a100, C4<1>, C4<1>;
v0x5c7c32e435f0_0 .net "in_a", 0 0, L_0x5c7c3311a100;  alias, 1 drivers
v0x5c7c32e436b0_0 .net "in_b", 0 0, L_0x5c7c3311a100;  alias, 1 drivers
v0x5c7c32e437a0_0 .net "out", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
S_0x5c7c32e43e50 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e41410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e44590_0 .net "in_a", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e44630_0 .net "out", 0 0, L_0x5c7c33119e40;  alias, 1 drivers
S_0x5c7c32e44020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e43e50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33119e40 .functor NAND 1, L_0x5c7c3311c320, L_0x5c7c3311c320, C4<1>, C4<1>;
v0x5c7c32e44270_0 .net "in_a", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e443c0_0 .net "in_b", 0 0, L_0x5c7c3311c320;  alias, 1 drivers
v0x5c7c32e44480_0 .net "out", 0 0, L_0x5c7c33119e40;  alias, 1 drivers
S_0x5c7c32e44730 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e41410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e44eb0_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e44f50_0 .net "out", 0 0, L_0x5c7c3311a050;  alias, 1 drivers
S_0x5c7c32e44950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e44730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a050 .functor NAND 1, L_0x5c7c3311c280, L_0x5c7c3311c280, C4<1>, C4<1>;
v0x5c7c32e44bc0_0 .net "in_a", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e44d10_0 .net "in_b", 0 0, L_0x5c7c3311c280;  alias, 1 drivers
v0x5c7c32e44dd0_0 .net "out", 0 0, L_0x5c7c3311a050;  alias, 1 drivers
S_0x5c7c32e45050 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e41410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e4ab20_0 .net "branch1_out", 0 0, L_0x5c7c3311a3c0;  1 drivers
v0x5c7c32e4ac50_0 .net "branch2_out", 0 0, L_0x5c7c3311a6e0;  1 drivers
v0x5c7c32e4ada0_0 .net "in_a", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
v0x5c7c32e4ae70_0 .net "in_b", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
v0x5c7c32e4af10_0 .net "out", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e4afb0_0 .net "temp1_out", 0 0, L_0x5c7c3311a310;  1 drivers
v0x5c7c32e4b050_0 .net "temp2_out", 0 0, L_0x5c7c3311a630;  1 drivers
v0x5c7c32e4b0f0_0 .net "temp3_out", 0 0, L_0x5c7c3311a950;  1 drivers
S_0x5c7c32e452d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e45050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e46360_0 .net "in_a", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
v0x5c7c32e46400_0 .net "in_b", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
v0x5c7c32e464c0_0 .net "out", 0 0, L_0x5c7c3311a310;  alias, 1 drivers
v0x5c7c32e465e0_0 .net "temp_out", 0 0, L_0x5c7c3311a260;  1 drivers
S_0x5c7c32e45540 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e452d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a260 .functor NAND 1, L_0x5c7c33119fa0, L_0x5c7c33119fa0, C4<1>, C4<1>;
v0x5c7c32e457b0_0 .net "in_a", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
v0x5c7c32e45870_0 .net "in_b", 0 0, L_0x5c7c33119fa0;  alias, 1 drivers
v0x5c7c32e459c0_0 .net "out", 0 0, L_0x5c7c3311a260;  alias, 1 drivers
S_0x5c7c32e45ac0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e452d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e461b0_0 .net "in_a", 0 0, L_0x5c7c3311a260;  alias, 1 drivers
v0x5c7c32e46250_0 .net "out", 0 0, L_0x5c7c3311a310;  alias, 1 drivers
S_0x5c7c32e45c90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e45ac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a310 .functor NAND 1, L_0x5c7c3311a260, L_0x5c7c3311a260, C4<1>, C4<1>;
v0x5c7c32e45f00_0 .net "in_a", 0 0, L_0x5c7c3311a260;  alias, 1 drivers
v0x5c7c32e45fc0_0 .net "in_b", 0 0, L_0x5c7c3311a260;  alias, 1 drivers
v0x5c7c32e460b0_0 .net "out", 0 0, L_0x5c7c3311a310;  alias, 1 drivers
S_0x5c7c32e46750 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e45050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e47780_0 .net "in_a", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
v0x5c7c32e47820_0 .net "in_b", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
v0x5c7c32e478e0_0 .net "out", 0 0, L_0x5c7c3311a630;  alias, 1 drivers
v0x5c7c32e47a00_0 .net "temp_out", 0 0, L_0x5c7c3311a580;  1 drivers
S_0x5c7c32e46930 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e46750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a580 .functor NAND 1, L_0x5c7c3311a1b0, L_0x5c7c3311a1b0, C4<1>, C4<1>;
v0x5c7c32e46ba0_0 .net "in_a", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
v0x5c7c32e46c60_0 .net "in_b", 0 0, L_0x5c7c3311a1b0;  alias, 1 drivers
v0x5c7c32e46db0_0 .net "out", 0 0, L_0x5c7c3311a580;  alias, 1 drivers
S_0x5c7c32e46eb0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e46750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e475d0_0 .net "in_a", 0 0, L_0x5c7c3311a580;  alias, 1 drivers
v0x5c7c32e47670_0 .net "out", 0 0, L_0x5c7c3311a630;  alias, 1 drivers
S_0x5c7c32e47080 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e46eb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a630 .functor NAND 1, L_0x5c7c3311a580, L_0x5c7c3311a580, C4<1>, C4<1>;
v0x5c7c32e472f0_0 .net "in_a", 0 0, L_0x5c7c3311a580;  alias, 1 drivers
v0x5c7c32e473e0_0 .net "in_b", 0 0, L_0x5c7c3311a580;  alias, 1 drivers
v0x5c7c32e474d0_0 .net "out", 0 0, L_0x5c7c3311a630;  alias, 1 drivers
S_0x5c7c32e47b70 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e45050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e48bb0_0 .net "in_a", 0 0, L_0x5c7c3311a3c0;  alias, 1 drivers
v0x5c7c32e48c80_0 .net "in_b", 0 0, L_0x5c7c3311a6e0;  alias, 1 drivers
v0x5c7c32e48d50_0 .net "out", 0 0, L_0x5c7c3311a950;  alias, 1 drivers
v0x5c7c32e48e70_0 .net "temp_out", 0 0, L_0x5c7c3311a8a0;  1 drivers
S_0x5c7c32e47d50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e47b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a8a0 .functor NAND 1, L_0x5c7c3311a3c0, L_0x5c7c3311a6e0, C4<1>, C4<1>;
v0x5c7c32e47fa0_0 .net "in_a", 0 0, L_0x5c7c3311a3c0;  alias, 1 drivers
v0x5c7c32e48080_0 .net "in_b", 0 0, L_0x5c7c3311a6e0;  alias, 1 drivers
v0x5c7c32e48140_0 .net "out", 0 0, L_0x5c7c3311a8a0;  alias, 1 drivers
S_0x5c7c32e48290 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e47b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e48a00_0 .net "in_a", 0 0, L_0x5c7c3311a8a0;  alias, 1 drivers
v0x5c7c32e48aa0_0 .net "out", 0 0, L_0x5c7c3311a950;  alias, 1 drivers
S_0x5c7c32e484b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e48290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a950 .functor NAND 1, L_0x5c7c3311a8a0, L_0x5c7c3311a8a0, C4<1>, C4<1>;
v0x5c7c32e48720_0 .net "in_a", 0 0, L_0x5c7c3311a8a0;  alias, 1 drivers
v0x5c7c32e48810_0 .net "in_b", 0 0, L_0x5c7c3311a8a0;  alias, 1 drivers
v0x5c7c32e48900_0 .net "out", 0 0, L_0x5c7c3311a950;  alias, 1 drivers
S_0x5c7c32e48fc0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e45050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e496f0_0 .net "in_a", 0 0, L_0x5c7c3311a310;  alias, 1 drivers
v0x5c7c32e49790_0 .net "out", 0 0, L_0x5c7c3311a3c0;  alias, 1 drivers
S_0x5c7c32e49190 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e48fc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a3c0 .functor NAND 1, L_0x5c7c3311a310, L_0x5c7c3311a310, C4<1>, C4<1>;
v0x5c7c32e49400_0 .net "in_a", 0 0, L_0x5c7c3311a310;  alias, 1 drivers
v0x5c7c32e494c0_0 .net "in_b", 0 0, L_0x5c7c3311a310;  alias, 1 drivers
v0x5c7c32e49610_0 .net "out", 0 0, L_0x5c7c3311a3c0;  alias, 1 drivers
S_0x5c7c32e49890 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e45050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e4a060_0 .net "in_a", 0 0, L_0x5c7c3311a630;  alias, 1 drivers
v0x5c7c32e4a100_0 .net "out", 0 0, L_0x5c7c3311a6e0;  alias, 1 drivers
S_0x5c7c32e49b00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e49890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311a6e0 .functor NAND 1, L_0x5c7c3311a630, L_0x5c7c3311a630, C4<1>, C4<1>;
v0x5c7c32e49d70_0 .net "in_a", 0 0, L_0x5c7c3311a630;  alias, 1 drivers
v0x5c7c32e49e30_0 .net "in_b", 0 0, L_0x5c7c3311a630;  alias, 1 drivers
v0x5c7c32e49f80_0 .net "out", 0 0, L_0x5c7c3311a6e0;  alias, 1 drivers
S_0x5c7c32e4a200 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e45050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e4a9a0_0 .net "in_a", 0 0, L_0x5c7c3311a950;  alias, 1 drivers
v0x5c7c32e4aa40_0 .net "out", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
S_0x5c7c32e4a420 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e4a200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311aa00 .functor NAND 1, L_0x5c7c3311a950, L_0x5c7c3311a950, C4<1>, C4<1>;
v0x5c7c32e4a690_0 .net "in_a", 0 0, L_0x5c7c3311a950;  alias, 1 drivers
v0x5c7c32e4a750_0 .net "in_b", 0 0, L_0x5c7c3311a950;  alias, 1 drivers
v0x5c7c32e4a8a0_0 .net "out", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
S_0x5c7c32e4bdb0 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32e3fad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e578d0_0 .net "a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e57970_0 .net "b", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e57a30_0 .net "carry", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e57ad0_0 .net "sum", 0 0, L_0x5c7c3311b930;  alias, 1 drivers
S_0x5c7c32e4bfd0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e4bdb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e4cf70_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e4d010_0 .net "in_b", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e4d0d0_0 .net "out", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e4d1f0_0 .net "temp_out", 0 0, L_0x5c7c32e4a830;  1 drivers
S_0x5c7c32e4c180 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e4bfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e4a830 .functor NAND 1, L_0x5c7c3311aa00, L_0x5c7c33119a20, C4<1>, C4<1>;
v0x5c7c32e4c3f0_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e4c4b0_0 .net "in_b", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e4c570_0 .net "out", 0 0, L_0x5c7c32e4a830;  alias, 1 drivers
S_0x5c7c32e4c6a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e4bfd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e4cdc0_0 .net "in_a", 0 0, L_0x5c7c32e4a830;  alias, 1 drivers
v0x5c7c32e4ce60_0 .net "out", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
S_0x5c7c32e4c870 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e4c6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b000 .functor NAND 1, L_0x5c7c32e4a830, L_0x5c7c32e4a830, C4<1>, C4<1>;
v0x5c7c32e4cae0_0 .net "in_a", 0 0, L_0x5c7c32e4a830;  alias, 1 drivers
v0x5c7c32e4cbd0_0 .net "in_b", 0 0, L_0x5c7c32e4a830;  alias, 1 drivers
v0x5c7c32e4ccc0_0 .net "out", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
S_0x5c7c32e4d360 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e4bdb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e571f0_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e57290_0 .net "in_b", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e57350_0 .net "out", 0 0, L_0x5c7c3311b930;  alias, 1 drivers
v0x5c7c32e573f0_0 .net "temp_a_and_out", 0 0, L_0x5c7c3311b210;  1 drivers
v0x5c7c32e575a0_0 .net "temp_a_out", 0 0, L_0x5c7c3311b0b0;  1 drivers
v0x5c7c32e57640_0 .net "temp_b_and_out", 0 0, L_0x5c7c3311b420;  1 drivers
v0x5c7c32e577f0_0 .net "temp_b_out", 0 0, L_0x5c7c3311b2c0;  1 drivers
S_0x5c7c32e4d540 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e4d360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e4e5e0_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e4e790_0 .net "in_b", 0 0, L_0x5c7c3311b0b0;  alias, 1 drivers
v0x5c7c32e4e880_0 .net "out", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
v0x5c7c32e4e9a0_0 .net "temp_out", 0 0, L_0x5c7c3311b160;  1 drivers
S_0x5c7c32e4d7b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e4d540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b160 .functor NAND 1, L_0x5c7c3311aa00, L_0x5c7c3311b0b0, C4<1>, C4<1>;
v0x5c7c32e4da20_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e4dae0_0 .net "in_b", 0 0, L_0x5c7c3311b0b0;  alias, 1 drivers
v0x5c7c32e4dba0_0 .net "out", 0 0, L_0x5c7c3311b160;  alias, 1 drivers
S_0x5c7c32e4dcc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e4d540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e4e430_0 .net "in_a", 0 0, L_0x5c7c3311b160;  alias, 1 drivers
v0x5c7c32e4e4d0_0 .net "out", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
S_0x5c7c32e4dee0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e4dcc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b210 .functor NAND 1, L_0x5c7c3311b160, L_0x5c7c3311b160, C4<1>, C4<1>;
v0x5c7c32e4e150_0 .net "in_a", 0 0, L_0x5c7c3311b160;  alias, 1 drivers
v0x5c7c32e4e240_0 .net "in_b", 0 0, L_0x5c7c3311b160;  alias, 1 drivers
v0x5c7c32e4e330_0 .net "out", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
S_0x5c7c32e4ea60 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e4d360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e4fa70_0 .net "in_a", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e4fb10_0 .net "in_b", 0 0, L_0x5c7c3311b2c0;  alias, 1 drivers
v0x5c7c32e4fc00_0 .net "out", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
v0x5c7c32e4fd20_0 .net "temp_out", 0 0, L_0x5c7c3311b370;  1 drivers
S_0x5c7c32e4ec40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e4ea60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b370 .functor NAND 1, L_0x5c7c33119a20, L_0x5c7c3311b2c0, C4<1>, C4<1>;
v0x5c7c32e4eeb0_0 .net "in_a", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e4ef70_0 .net "in_b", 0 0, L_0x5c7c3311b2c0;  alias, 1 drivers
v0x5c7c32e4f030_0 .net "out", 0 0, L_0x5c7c3311b370;  alias, 1 drivers
S_0x5c7c32e4f150 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e4ea60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e4f8c0_0 .net "in_a", 0 0, L_0x5c7c3311b370;  alias, 1 drivers
v0x5c7c32e4f960_0 .net "out", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
S_0x5c7c32e4f370 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e4f150;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b420 .functor NAND 1, L_0x5c7c3311b370, L_0x5c7c3311b370, C4<1>, C4<1>;
v0x5c7c32e4f5e0_0 .net "in_a", 0 0, L_0x5c7c3311b370;  alias, 1 drivers
v0x5c7c32e4f6d0_0 .net "in_b", 0 0, L_0x5c7c3311b370;  alias, 1 drivers
v0x5c7c32e4f7c0_0 .net "out", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
S_0x5c7c32e4fe70 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e4d360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e50680_0 .net "in_a", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e50720_0 .net "out", 0 0, L_0x5c7c3311b0b0;  alias, 1 drivers
S_0x5c7c32e50040 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e4fe70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b0b0 .functor NAND 1, L_0x5c7c33119a20, L_0x5c7c33119a20, C4<1>, C4<1>;
v0x5c7c32e50290_0 .net "in_a", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e50460_0 .net "in_b", 0 0, L_0x5c7c33119a20;  alias, 1 drivers
v0x5c7c32e50520_0 .net "out", 0 0, L_0x5c7c3311b0b0;  alias, 1 drivers
S_0x5c7c32e50820 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e4d360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e50f60_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e51000_0 .net "out", 0 0, L_0x5c7c3311b2c0;  alias, 1 drivers
S_0x5c7c32e50a40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e50820;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b2c0 .functor NAND 1, L_0x5c7c3311aa00, L_0x5c7c3311aa00, C4<1>, C4<1>;
v0x5c7c32e50cb0_0 .net "in_a", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e50d70_0 .net "in_b", 0 0, L_0x5c7c3311aa00;  alias, 1 drivers
v0x5c7c32e50e30_0 .net "out", 0 0, L_0x5c7c3311b2c0;  alias, 1 drivers
S_0x5c7c32e51100 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e4d360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e56b40_0 .net "branch1_out", 0 0, L_0x5c7c3311b630;  1 drivers
v0x5c7c32e56c70_0 .net "branch2_out", 0 0, L_0x5c7c3311b7b0;  1 drivers
v0x5c7c32e56dc0_0 .net "in_a", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
v0x5c7c32e56e90_0 .net "in_b", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
v0x5c7c32e56f30_0 .net "out", 0 0, L_0x5c7c3311b930;  alias, 1 drivers
v0x5c7c32e56fd0_0 .net "temp1_out", 0 0, L_0x5c7c3311b580;  1 drivers
v0x5c7c32e57070_0 .net "temp2_out", 0 0, L_0x5c7c3311b700;  1 drivers
v0x5c7c32e57110_0 .net "temp3_out", 0 0, L_0x5c7c3311b880;  1 drivers
S_0x5c7c32e51380 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e51100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e52380_0 .net "in_a", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
v0x5c7c32e52420_0 .net "in_b", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
v0x5c7c32e524e0_0 .net "out", 0 0, L_0x5c7c3311b580;  alias, 1 drivers
v0x5c7c32e52600_0 .net "temp_out", 0 0, L_0x5c7c3311b4d0;  1 drivers
S_0x5c7c32e515f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e51380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b4d0 .functor NAND 1, L_0x5c7c3311b210, L_0x5c7c3311b210, C4<1>, C4<1>;
v0x5c7c32e51860_0 .net "in_a", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
v0x5c7c32e51920_0 .net "in_b", 0 0, L_0x5c7c3311b210;  alias, 1 drivers
v0x5c7c32e519e0_0 .net "out", 0 0, L_0x5c7c3311b4d0;  alias, 1 drivers
S_0x5c7c32e51ae0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e51380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e521d0_0 .net "in_a", 0 0, L_0x5c7c3311b4d0;  alias, 1 drivers
v0x5c7c32e52270_0 .net "out", 0 0, L_0x5c7c3311b580;  alias, 1 drivers
S_0x5c7c32e51cb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e51ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b580 .functor NAND 1, L_0x5c7c3311b4d0, L_0x5c7c3311b4d0, C4<1>, C4<1>;
v0x5c7c32e51f20_0 .net "in_a", 0 0, L_0x5c7c3311b4d0;  alias, 1 drivers
v0x5c7c32e51fe0_0 .net "in_b", 0 0, L_0x5c7c3311b4d0;  alias, 1 drivers
v0x5c7c32e520d0_0 .net "out", 0 0, L_0x5c7c3311b580;  alias, 1 drivers
S_0x5c7c32e52770 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e51100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e537a0_0 .net "in_a", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
v0x5c7c32e53840_0 .net "in_b", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
v0x5c7c32e53900_0 .net "out", 0 0, L_0x5c7c3311b700;  alias, 1 drivers
v0x5c7c32e53a20_0 .net "temp_out", 0 0, L_0x5c7c32e555c0;  1 drivers
S_0x5c7c32e52950 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e52770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e555c0 .functor NAND 1, L_0x5c7c3311b420, L_0x5c7c3311b420, C4<1>, C4<1>;
v0x5c7c32e52bc0_0 .net "in_a", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
v0x5c7c32e52c80_0 .net "in_b", 0 0, L_0x5c7c3311b420;  alias, 1 drivers
v0x5c7c32e52dd0_0 .net "out", 0 0, L_0x5c7c32e555c0;  alias, 1 drivers
S_0x5c7c32e52ed0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e52770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e535f0_0 .net "in_a", 0 0, L_0x5c7c32e555c0;  alias, 1 drivers
v0x5c7c32e53690_0 .net "out", 0 0, L_0x5c7c3311b700;  alias, 1 drivers
S_0x5c7c32e530a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e52ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b700 .functor NAND 1, L_0x5c7c32e555c0, L_0x5c7c32e555c0, C4<1>, C4<1>;
v0x5c7c32e53310_0 .net "in_a", 0 0, L_0x5c7c32e555c0;  alias, 1 drivers
v0x5c7c32e53400_0 .net "in_b", 0 0, L_0x5c7c32e555c0;  alias, 1 drivers
v0x5c7c32e534f0_0 .net "out", 0 0, L_0x5c7c3311b700;  alias, 1 drivers
S_0x5c7c32e53b90 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e51100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e54bd0_0 .net "in_a", 0 0, L_0x5c7c3311b630;  alias, 1 drivers
v0x5c7c32e54ca0_0 .net "in_b", 0 0, L_0x5c7c3311b7b0;  alias, 1 drivers
v0x5c7c32e54d70_0 .net "out", 0 0, L_0x5c7c3311b880;  alias, 1 drivers
v0x5c7c32e54e90_0 .net "temp_out", 0 0, L_0x5c7c32e55f30;  1 drivers
S_0x5c7c32e53d70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e53b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e55f30 .functor NAND 1, L_0x5c7c3311b630, L_0x5c7c3311b7b0, C4<1>, C4<1>;
v0x5c7c32e53fc0_0 .net "in_a", 0 0, L_0x5c7c3311b630;  alias, 1 drivers
v0x5c7c32e540a0_0 .net "in_b", 0 0, L_0x5c7c3311b7b0;  alias, 1 drivers
v0x5c7c32e54160_0 .net "out", 0 0, L_0x5c7c32e55f30;  alias, 1 drivers
S_0x5c7c32e542b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e53b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e54a20_0 .net "in_a", 0 0, L_0x5c7c32e55f30;  alias, 1 drivers
v0x5c7c32e54ac0_0 .net "out", 0 0, L_0x5c7c3311b880;  alias, 1 drivers
S_0x5c7c32e544d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e542b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b880 .functor NAND 1, L_0x5c7c32e55f30, L_0x5c7c32e55f30, C4<1>, C4<1>;
v0x5c7c32e54740_0 .net "in_a", 0 0, L_0x5c7c32e55f30;  alias, 1 drivers
v0x5c7c32e54830_0 .net "in_b", 0 0, L_0x5c7c32e55f30;  alias, 1 drivers
v0x5c7c32e54920_0 .net "out", 0 0, L_0x5c7c3311b880;  alias, 1 drivers
S_0x5c7c32e54fe0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e51100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e55710_0 .net "in_a", 0 0, L_0x5c7c3311b580;  alias, 1 drivers
v0x5c7c32e557b0_0 .net "out", 0 0, L_0x5c7c3311b630;  alias, 1 drivers
S_0x5c7c32e551b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e54fe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b630 .functor NAND 1, L_0x5c7c3311b580, L_0x5c7c3311b580, C4<1>, C4<1>;
v0x5c7c32e55420_0 .net "in_a", 0 0, L_0x5c7c3311b580;  alias, 1 drivers
v0x5c7c32e554e0_0 .net "in_b", 0 0, L_0x5c7c3311b580;  alias, 1 drivers
v0x5c7c32e55630_0 .net "out", 0 0, L_0x5c7c3311b630;  alias, 1 drivers
S_0x5c7c32e558b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e51100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e56080_0 .net "in_a", 0 0, L_0x5c7c3311b700;  alias, 1 drivers
v0x5c7c32e56120_0 .net "out", 0 0, L_0x5c7c3311b7b0;  alias, 1 drivers
S_0x5c7c32e55b20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e558b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b7b0 .functor NAND 1, L_0x5c7c3311b700, L_0x5c7c3311b700, C4<1>, C4<1>;
v0x5c7c32e55d90_0 .net "in_a", 0 0, L_0x5c7c3311b700;  alias, 1 drivers
v0x5c7c32e55e50_0 .net "in_b", 0 0, L_0x5c7c3311b700;  alias, 1 drivers
v0x5c7c32e55fa0_0 .net "out", 0 0, L_0x5c7c3311b7b0;  alias, 1 drivers
S_0x5c7c32e56220 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e51100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e569c0_0 .net "in_a", 0 0, L_0x5c7c3311b880;  alias, 1 drivers
v0x5c7c32e56a60_0 .net "out", 0 0, L_0x5c7c3311b930;  alias, 1 drivers
S_0x5c7c32e56440 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e56220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311b930 .functor NAND 1, L_0x5c7c3311b880, L_0x5c7c3311b880, C4<1>, C4<1>;
v0x5c7c32e566b0_0 .net "in_a", 0 0, L_0x5c7c3311b880;  alias, 1 drivers
v0x5c7c32e56770_0 .net "in_b", 0 0, L_0x5c7c3311b880;  alias, 1 drivers
v0x5c7c32e568c0_0 .net "out", 0 0, L_0x5c7c3311b930;  alias, 1 drivers
S_0x5c7c32e57c40 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32e3fad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e5d630_0 .net "branch1_out", 0 0, L_0x5c7c3311bbc0;  1 drivers
v0x5c7c32e5d760_0 .net "branch2_out", 0 0, L_0x5c7c3311be50;  1 drivers
v0x5c7c32e5d8b0_0 .net "in_a", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e5da90_0 .net "in_b", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e5dc40_0 .net "out", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e5dce0_0 .net "temp1_out", 0 0, L_0x5c7c3311bb10;  1 drivers
v0x5c7c32e5dd80_0 .net "temp2_out", 0 0, L_0x5c7c3311bda0;  1 drivers
v0x5c7c32e5de20_0 .net "temp3_out", 0 0, L_0x5c7c3311c030;  1 drivers
S_0x5c7c32e57dd0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e57c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e58e70_0 .net "in_a", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e58f10_0 .net "in_b", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e58fd0_0 .net "out", 0 0, L_0x5c7c3311bb10;  alias, 1 drivers
v0x5c7c32e590f0_0 .net "temp_out", 0 0, L_0x5c7c32e56850;  1 drivers
S_0x5c7c32e57ff0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e57dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e56850 .functor NAND 1, L_0x5c7c33119d90, L_0x5c7c33119d90, C4<1>, C4<1>;
v0x5c7c32e58260_0 .net "in_a", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e583b0_0 .net "in_b", 0 0, L_0x5c7c33119d90;  alias, 1 drivers
v0x5c7c32e58470_0 .net "out", 0 0, L_0x5c7c32e56850;  alias, 1 drivers
S_0x5c7c32e585a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e57dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e58cc0_0 .net "in_a", 0 0, L_0x5c7c32e56850;  alias, 1 drivers
v0x5c7c32e58d60_0 .net "out", 0 0, L_0x5c7c3311bb10;  alias, 1 drivers
S_0x5c7c32e58770 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e585a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311bb10 .functor NAND 1, L_0x5c7c32e56850, L_0x5c7c32e56850, C4<1>, C4<1>;
v0x5c7c32e589e0_0 .net "in_a", 0 0, L_0x5c7c32e56850;  alias, 1 drivers
v0x5c7c32e58ad0_0 .net "in_b", 0 0, L_0x5c7c32e56850;  alias, 1 drivers
v0x5c7c32e58bc0_0 .net "out", 0 0, L_0x5c7c3311bb10;  alias, 1 drivers
S_0x5c7c32e59260 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e57c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e5a290_0 .net "in_a", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e5a330_0 .net "in_b", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e5a3f0_0 .net "out", 0 0, L_0x5c7c3311bda0;  alias, 1 drivers
v0x5c7c32e5a510_0 .net "temp_out", 0 0, L_0x5c7c32e5c0b0;  1 drivers
S_0x5c7c32e59440 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e59260;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e5c0b0 .functor NAND 1, L_0x5c7c3311b000, L_0x5c7c3311b000, C4<1>, C4<1>;
v0x5c7c32e596b0_0 .net "in_a", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e59800_0 .net "in_b", 0 0, L_0x5c7c3311b000;  alias, 1 drivers
v0x5c7c32e598c0_0 .net "out", 0 0, L_0x5c7c32e5c0b0;  alias, 1 drivers
S_0x5c7c32e599c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e59260;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e5a0e0_0 .net "in_a", 0 0, L_0x5c7c32e5c0b0;  alias, 1 drivers
v0x5c7c32e5a180_0 .net "out", 0 0, L_0x5c7c3311bda0;  alias, 1 drivers
S_0x5c7c32e59b90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e599c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311bda0 .functor NAND 1, L_0x5c7c32e5c0b0, L_0x5c7c32e5c0b0, C4<1>, C4<1>;
v0x5c7c32e59e00_0 .net "in_a", 0 0, L_0x5c7c32e5c0b0;  alias, 1 drivers
v0x5c7c32e59ef0_0 .net "in_b", 0 0, L_0x5c7c32e5c0b0;  alias, 1 drivers
v0x5c7c32e59fe0_0 .net "out", 0 0, L_0x5c7c3311bda0;  alias, 1 drivers
S_0x5c7c32e5a680 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e57c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e5b6c0_0 .net "in_a", 0 0, L_0x5c7c3311bbc0;  alias, 1 drivers
v0x5c7c32e5b790_0 .net "in_b", 0 0, L_0x5c7c3311be50;  alias, 1 drivers
v0x5c7c32e5b860_0 .net "out", 0 0, L_0x5c7c3311c030;  alias, 1 drivers
v0x5c7c32e5b980_0 .net "temp_out", 0 0, L_0x5c7c32e5ca20;  1 drivers
S_0x5c7c32e5a860 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e5a680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e5ca20 .functor NAND 1, L_0x5c7c3311bbc0, L_0x5c7c3311be50, C4<1>, C4<1>;
v0x5c7c32e5aab0_0 .net "in_a", 0 0, L_0x5c7c3311bbc0;  alias, 1 drivers
v0x5c7c32e5ab90_0 .net "in_b", 0 0, L_0x5c7c3311be50;  alias, 1 drivers
v0x5c7c32e5ac50_0 .net "out", 0 0, L_0x5c7c32e5ca20;  alias, 1 drivers
S_0x5c7c32e5ada0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e5a680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e5b510_0 .net "in_a", 0 0, L_0x5c7c32e5ca20;  alias, 1 drivers
v0x5c7c32e5b5b0_0 .net "out", 0 0, L_0x5c7c3311c030;  alias, 1 drivers
S_0x5c7c32e5afc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e5ada0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c030 .functor NAND 1, L_0x5c7c32e5ca20, L_0x5c7c32e5ca20, C4<1>, C4<1>;
v0x5c7c32e5b230_0 .net "in_a", 0 0, L_0x5c7c32e5ca20;  alias, 1 drivers
v0x5c7c32e5b320_0 .net "in_b", 0 0, L_0x5c7c32e5ca20;  alias, 1 drivers
v0x5c7c32e5b410_0 .net "out", 0 0, L_0x5c7c3311c030;  alias, 1 drivers
S_0x5c7c32e5bad0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e57c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e5c200_0 .net "in_a", 0 0, L_0x5c7c3311bb10;  alias, 1 drivers
v0x5c7c32e5c2a0_0 .net "out", 0 0, L_0x5c7c3311bbc0;  alias, 1 drivers
S_0x5c7c32e5bca0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e5bad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311bbc0 .functor NAND 1, L_0x5c7c3311bb10, L_0x5c7c3311bb10, C4<1>, C4<1>;
v0x5c7c32e5bf10_0 .net "in_a", 0 0, L_0x5c7c3311bb10;  alias, 1 drivers
v0x5c7c32e5bfd0_0 .net "in_b", 0 0, L_0x5c7c3311bb10;  alias, 1 drivers
v0x5c7c32e5c120_0 .net "out", 0 0, L_0x5c7c3311bbc0;  alias, 1 drivers
S_0x5c7c32e5c3a0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e57c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e5cb70_0 .net "in_a", 0 0, L_0x5c7c3311bda0;  alias, 1 drivers
v0x5c7c32e5cc10_0 .net "out", 0 0, L_0x5c7c3311be50;  alias, 1 drivers
S_0x5c7c32e5c610 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e5c3a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311be50 .functor NAND 1, L_0x5c7c3311bda0, L_0x5c7c3311bda0, C4<1>, C4<1>;
v0x5c7c32e5c880_0 .net "in_a", 0 0, L_0x5c7c3311bda0;  alias, 1 drivers
v0x5c7c32e5c940_0 .net "in_b", 0 0, L_0x5c7c3311bda0;  alias, 1 drivers
v0x5c7c32e5ca90_0 .net "out", 0 0, L_0x5c7c3311be50;  alias, 1 drivers
S_0x5c7c32e5cd10 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e57c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e5d4b0_0 .net "in_a", 0 0, L_0x5c7c3311c030;  alias, 1 drivers
v0x5c7c32e5d550_0 .net "out", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
S_0x5c7c32e5cf30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e5cd10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c0e0 .functor NAND 1, L_0x5c7c3311c030, L_0x5c7c3311c030, C4<1>, C4<1>;
v0x5c7c32e5d1a0_0 .net "in_a", 0 0, L_0x5c7c3311c030;  alias, 1 drivers
v0x5c7c32e5d260_0 .net "in_b", 0 0, L_0x5c7c3311c030;  alias, 1 drivers
v0x5c7c32e5d3b0_0 .net "out", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
S_0x5c7c32e5e480 .scope module, "fa_gate6" "FullAdder" 2 11, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32e7c8b0_0 .net "a", 0 0, L_0x5c7c3311e840;  1 drivers
v0x5c7c32e7c950_0 .net "b", 0 0, L_0x5c7c3311e8e0;  1 drivers
v0x5c7c32e7ca10_0 .net "c", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e7cab0_0 .net "carry", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e7cb50_0 .net "sum", 0 0, L_0x5c7c3311def0;  1 drivers
v0x5c7c32e7cbf0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c3311c470;  1 drivers
v0x5c7c32e7cc90_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c3311d5c0;  1 drivers
v0x5c7c32e7cd30_0 .net "tmp_sum_out", 0 0, L_0x5c7c3311cfc0;  1 drivers
S_0x5c7c32e5e6e0 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32e5e480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e6a260_0 .net "a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e6a410_0 .net "b", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e6a5e0_0 .net "carry", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e6a680_0 .net "sum", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
S_0x5c7c32e5e950 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e5e6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e5fa40_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e5fb10_0 .net "in_b", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e5fbe0_0 .net "out", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e5fd00_0 .net "temp_out", 0 0, L_0x5c7c3311c3c0;  1 drivers
S_0x5c7c32e5ebc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e5e950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c3c0 .functor NAND 1, L_0x5c7c3311e840, L_0x5c7c3311e8e0, C4<1>, C4<1>;
v0x5c7c32e5ee30_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e5ef10_0 .net "in_b", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e5efd0_0 .net "out", 0 0, L_0x5c7c3311c3c0;  alias, 1 drivers
S_0x5c7c32e5f120 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e5e950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e5f890_0 .net "in_a", 0 0, L_0x5c7c3311c3c0;  alias, 1 drivers
v0x5c7c32e5f930_0 .net "out", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
S_0x5c7c32e5f340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e5f120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c470 .functor NAND 1, L_0x5c7c3311c3c0, L_0x5c7c3311c3c0, C4<1>, C4<1>;
v0x5c7c32e5f5b0_0 .net "in_a", 0 0, L_0x5c7c3311c3c0;  alias, 1 drivers
v0x5c7c32e5f6a0_0 .net "in_b", 0 0, L_0x5c7c3311c3c0;  alias, 1 drivers
v0x5c7c32e5f790_0 .net "out", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
S_0x5c7c32e5fdc0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e5e6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e69b80_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e69c20_0 .net "in_b", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e69ce0_0 .net "out", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e69d80_0 .net "temp_a_and_out", 0 0, L_0x5c7c3311c680;  1 drivers
v0x5c7c32e69f30_0 .net "temp_a_out", 0 0, L_0x5c7c3311c520;  1 drivers
v0x5c7c32e69fd0_0 .net "temp_b_and_out", 0 0, L_0x5c7c3311c890;  1 drivers
v0x5c7c32e6a180_0 .net "temp_b_out", 0 0, L_0x5c7c3311c730;  1 drivers
S_0x5c7c32e5ffa0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e5fdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e61060_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e61100_0 .net "in_b", 0 0, L_0x5c7c3311c520;  alias, 1 drivers
v0x5c7c32e611f0_0 .net "out", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
v0x5c7c32e61310_0 .net "temp_out", 0 0, L_0x5c7c3311c5d0;  1 drivers
S_0x5c7c32e60210 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e5ffa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c5d0 .functor NAND 1, L_0x5c7c3311e840, L_0x5c7c3311c520, C4<1>, C4<1>;
v0x5c7c32e60480_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e60590_0 .net "in_b", 0 0, L_0x5c7c3311c520;  alias, 1 drivers
v0x5c7c32e60650_0 .net "out", 0 0, L_0x5c7c3311c5d0;  alias, 1 drivers
S_0x5c7c32e60770 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e5ffa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e60eb0_0 .net "in_a", 0 0, L_0x5c7c3311c5d0;  alias, 1 drivers
v0x5c7c32e60f50_0 .net "out", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
S_0x5c7c32e60990 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e60770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c680 .functor NAND 1, L_0x5c7c3311c5d0, L_0x5c7c3311c5d0, C4<1>, C4<1>;
v0x5c7c32e60c00_0 .net "in_a", 0 0, L_0x5c7c3311c5d0;  alias, 1 drivers
v0x5c7c32e60cc0_0 .net "in_b", 0 0, L_0x5c7c3311c5d0;  alias, 1 drivers
v0x5c7c32e60db0_0 .net "out", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
S_0x5c7c32e613d0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e5fdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e62400_0 .net "in_a", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e624a0_0 .net "in_b", 0 0, L_0x5c7c3311c730;  alias, 1 drivers
v0x5c7c32e62590_0 .net "out", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
v0x5c7c32e626b0_0 .net "temp_out", 0 0, L_0x5c7c3311c7e0;  1 drivers
S_0x5c7c32e615b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e613d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c7e0 .functor NAND 1, L_0x5c7c3311e8e0, L_0x5c7c3311c730, C4<1>, C4<1>;
v0x5c7c32e61820_0 .net "in_a", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e61930_0 .net "in_b", 0 0, L_0x5c7c3311c730;  alias, 1 drivers
v0x5c7c32e619f0_0 .net "out", 0 0, L_0x5c7c3311c7e0;  alias, 1 drivers
S_0x5c7c32e61b10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e613d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e62250_0 .net "in_a", 0 0, L_0x5c7c3311c7e0;  alias, 1 drivers
v0x5c7c32e622f0_0 .net "out", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
S_0x5c7c32e61d30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e61b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c890 .functor NAND 1, L_0x5c7c3311c7e0, L_0x5c7c3311c7e0, C4<1>, C4<1>;
v0x5c7c32e61fa0_0 .net "in_a", 0 0, L_0x5c7c3311c7e0;  alias, 1 drivers
v0x5c7c32e62060_0 .net "in_b", 0 0, L_0x5c7c3311c7e0;  alias, 1 drivers
v0x5c7c32e62150_0 .net "out", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
S_0x5c7c32e62800 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e5fdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e62f40_0 .net "in_a", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e62fe0_0 .net "out", 0 0, L_0x5c7c3311c520;  alias, 1 drivers
S_0x5c7c32e629d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e62800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c520 .functor NAND 1, L_0x5c7c3311e8e0, L_0x5c7c3311e8e0, C4<1>, C4<1>;
v0x5c7c32e62c20_0 .net "in_a", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e62d70_0 .net "in_b", 0 0, L_0x5c7c3311e8e0;  alias, 1 drivers
v0x5c7c32e62e30_0 .net "out", 0 0, L_0x5c7c3311c520;  alias, 1 drivers
S_0x5c7c32e630e0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e5fdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e63860_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e63900_0 .net "out", 0 0, L_0x5c7c3311c730;  alias, 1 drivers
S_0x5c7c32e63300 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e630e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c730 .functor NAND 1, L_0x5c7c3311e840, L_0x5c7c3311e840, C4<1>, C4<1>;
v0x5c7c32e63570_0 .net "in_a", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e636c0_0 .net "in_b", 0 0, L_0x5c7c3311e840;  alias, 1 drivers
v0x5c7c32e63780_0 .net "out", 0 0, L_0x5c7c3311c730;  alias, 1 drivers
S_0x5c7c32e63a00 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e5fdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e694d0_0 .net "branch1_out", 0 0, L_0x5c7c3311caa0;  1 drivers
v0x5c7c32e69600_0 .net "branch2_out", 0 0, L_0x5c7c3311cd30;  1 drivers
v0x5c7c32e69750_0 .net "in_a", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
v0x5c7c32e69820_0 .net "in_b", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
v0x5c7c32e698c0_0 .net "out", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e69960_0 .net "temp1_out", 0 0, L_0x5c7c3311c9f0;  1 drivers
v0x5c7c32e69a00_0 .net "temp2_out", 0 0, L_0x5c7c3311cc80;  1 drivers
v0x5c7c32e69aa0_0 .net "temp3_out", 0 0, L_0x5c7c3311cf10;  1 drivers
S_0x5c7c32e63c80 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e63a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e64d10_0 .net "in_a", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
v0x5c7c32e64db0_0 .net "in_b", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
v0x5c7c32e64e70_0 .net "out", 0 0, L_0x5c7c3311c9f0;  alias, 1 drivers
v0x5c7c32e64f90_0 .net "temp_out", 0 0, L_0x5c7c3311c940;  1 drivers
S_0x5c7c32e63ef0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e63c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c940 .functor NAND 1, L_0x5c7c3311c680, L_0x5c7c3311c680, C4<1>, C4<1>;
v0x5c7c32e64160_0 .net "in_a", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
v0x5c7c32e64220_0 .net "in_b", 0 0, L_0x5c7c3311c680;  alias, 1 drivers
v0x5c7c32e64370_0 .net "out", 0 0, L_0x5c7c3311c940;  alias, 1 drivers
S_0x5c7c32e64470 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e63c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e64b60_0 .net "in_a", 0 0, L_0x5c7c3311c940;  alias, 1 drivers
v0x5c7c32e64c00_0 .net "out", 0 0, L_0x5c7c3311c9f0;  alias, 1 drivers
S_0x5c7c32e64640 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e64470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311c9f0 .functor NAND 1, L_0x5c7c3311c940, L_0x5c7c3311c940, C4<1>, C4<1>;
v0x5c7c32e648b0_0 .net "in_a", 0 0, L_0x5c7c3311c940;  alias, 1 drivers
v0x5c7c32e64970_0 .net "in_b", 0 0, L_0x5c7c3311c940;  alias, 1 drivers
v0x5c7c32e64a60_0 .net "out", 0 0, L_0x5c7c3311c9f0;  alias, 1 drivers
S_0x5c7c32e65100 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e63a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e66130_0 .net "in_a", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
v0x5c7c32e661d0_0 .net "in_b", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
v0x5c7c32e66290_0 .net "out", 0 0, L_0x5c7c3311cc80;  alias, 1 drivers
v0x5c7c32e663b0_0 .net "temp_out", 0 0, L_0x5c7c32e67f50;  1 drivers
S_0x5c7c32e652e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e65100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e67f50 .functor NAND 1, L_0x5c7c3311c890, L_0x5c7c3311c890, C4<1>, C4<1>;
v0x5c7c32e65550_0 .net "in_a", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
v0x5c7c32e65610_0 .net "in_b", 0 0, L_0x5c7c3311c890;  alias, 1 drivers
v0x5c7c32e65760_0 .net "out", 0 0, L_0x5c7c32e67f50;  alias, 1 drivers
S_0x5c7c32e65860 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e65100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e65f80_0 .net "in_a", 0 0, L_0x5c7c32e67f50;  alias, 1 drivers
v0x5c7c32e66020_0 .net "out", 0 0, L_0x5c7c3311cc80;  alias, 1 drivers
S_0x5c7c32e65a30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e65860;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311cc80 .functor NAND 1, L_0x5c7c32e67f50, L_0x5c7c32e67f50, C4<1>, C4<1>;
v0x5c7c32e65ca0_0 .net "in_a", 0 0, L_0x5c7c32e67f50;  alias, 1 drivers
v0x5c7c32e65d90_0 .net "in_b", 0 0, L_0x5c7c32e67f50;  alias, 1 drivers
v0x5c7c32e65e80_0 .net "out", 0 0, L_0x5c7c3311cc80;  alias, 1 drivers
S_0x5c7c32e66520 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e63a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e67560_0 .net "in_a", 0 0, L_0x5c7c3311caa0;  alias, 1 drivers
v0x5c7c32e67630_0 .net "in_b", 0 0, L_0x5c7c3311cd30;  alias, 1 drivers
v0x5c7c32e67700_0 .net "out", 0 0, L_0x5c7c3311cf10;  alias, 1 drivers
v0x5c7c32e67820_0 .net "temp_out", 0 0, L_0x5c7c32e688c0;  1 drivers
S_0x5c7c32e66700 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e66520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e688c0 .functor NAND 1, L_0x5c7c3311caa0, L_0x5c7c3311cd30, C4<1>, C4<1>;
v0x5c7c32e66950_0 .net "in_a", 0 0, L_0x5c7c3311caa0;  alias, 1 drivers
v0x5c7c32e66a30_0 .net "in_b", 0 0, L_0x5c7c3311cd30;  alias, 1 drivers
v0x5c7c32e66af0_0 .net "out", 0 0, L_0x5c7c32e688c0;  alias, 1 drivers
S_0x5c7c32e66c40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e66520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e673b0_0 .net "in_a", 0 0, L_0x5c7c32e688c0;  alias, 1 drivers
v0x5c7c32e67450_0 .net "out", 0 0, L_0x5c7c3311cf10;  alias, 1 drivers
S_0x5c7c32e66e60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e66c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311cf10 .functor NAND 1, L_0x5c7c32e688c0, L_0x5c7c32e688c0, C4<1>, C4<1>;
v0x5c7c32e670d0_0 .net "in_a", 0 0, L_0x5c7c32e688c0;  alias, 1 drivers
v0x5c7c32e671c0_0 .net "in_b", 0 0, L_0x5c7c32e688c0;  alias, 1 drivers
v0x5c7c32e672b0_0 .net "out", 0 0, L_0x5c7c3311cf10;  alias, 1 drivers
S_0x5c7c32e67970 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e63a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e680a0_0 .net "in_a", 0 0, L_0x5c7c3311c9f0;  alias, 1 drivers
v0x5c7c32e68140_0 .net "out", 0 0, L_0x5c7c3311caa0;  alias, 1 drivers
S_0x5c7c32e67b40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e67970;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311caa0 .functor NAND 1, L_0x5c7c3311c9f0, L_0x5c7c3311c9f0, C4<1>, C4<1>;
v0x5c7c32e67db0_0 .net "in_a", 0 0, L_0x5c7c3311c9f0;  alias, 1 drivers
v0x5c7c32e67e70_0 .net "in_b", 0 0, L_0x5c7c3311c9f0;  alias, 1 drivers
v0x5c7c32e67fc0_0 .net "out", 0 0, L_0x5c7c3311caa0;  alias, 1 drivers
S_0x5c7c32e68240 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e63a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e68a10_0 .net "in_a", 0 0, L_0x5c7c3311cc80;  alias, 1 drivers
v0x5c7c32e68ab0_0 .net "out", 0 0, L_0x5c7c3311cd30;  alias, 1 drivers
S_0x5c7c32e684b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e68240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311cd30 .functor NAND 1, L_0x5c7c3311cc80, L_0x5c7c3311cc80, C4<1>, C4<1>;
v0x5c7c32e68720_0 .net "in_a", 0 0, L_0x5c7c3311cc80;  alias, 1 drivers
v0x5c7c32e687e0_0 .net "in_b", 0 0, L_0x5c7c3311cc80;  alias, 1 drivers
v0x5c7c32e68930_0 .net "out", 0 0, L_0x5c7c3311cd30;  alias, 1 drivers
S_0x5c7c32e68bb0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e63a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e69350_0 .net "in_a", 0 0, L_0x5c7c3311cf10;  alias, 1 drivers
v0x5c7c32e693f0_0 .net "out", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
S_0x5c7c32e68dd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e68bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311cfc0 .functor NAND 1, L_0x5c7c3311cf10, L_0x5c7c3311cf10, C4<1>, C4<1>;
v0x5c7c32e69040_0 .net "in_a", 0 0, L_0x5c7c3311cf10;  alias, 1 drivers
v0x5c7c32e69100_0 .net "in_b", 0 0, L_0x5c7c3311cf10;  alias, 1 drivers
v0x5c7c32e69250_0 .net "out", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
S_0x5c7c32e6a760 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32e5e480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e76280_0 .net "a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e76320_0 .net "b", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e763e0_0 .net "carry", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e76480_0 .net "sum", 0 0, L_0x5c7c3311def0;  alias, 1 drivers
S_0x5c7c32e6a980 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e6a760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e6b920_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6b9c0_0 .net "in_b", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6ba80_0 .net "out", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e6bba0_0 .net "temp_out", 0 0, L_0x5c7c32e691e0;  1 drivers
S_0x5c7c32e6ab30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e6a980;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e691e0 .functor NAND 1, L_0x5c7c3311cfc0, L_0x5c7c3311c0e0, C4<1>, C4<1>;
v0x5c7c32e6ada0_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6ae60_0 .net "in_b", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6af20_0 .net "out", 0 0, L_0x5c7c32e691e0;  alias, 1 drivers
S_0x5c7c32e6b050 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e6a980;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e6b770_0 .net "in_a", 0 0, L_0x5c7c32e691e0;  alias, 1 drivers
v0x5c7c32e6b810_0 .net "out", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
S_0x5c7c32e6b220 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e6b050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d5c0 .functor NAND 1, L_0x5c7c32e691e0, L_0x5c7c32e691e0, C4<1>, C4<1>;
v0x5c7c32e6b490_0 .net "in_a", 0 0, L_0x5c7c32e691e0;  alias, 1 drivers
v0x5c7c32e6b580_0 .net "in_b", 0 0, L_0x5c7c32e691e0;  alias, 1 drivers
v0x5c7c32e6b670_0 .net "out", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
S_0x5c7c32e6bd10 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e6a760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e75ba0_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e75c40_0 .net "in_b", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e75d00_0 .net "out", 0 0, L_0x5c7c3311def0;  alias, 1 drivers
v0x5c7c32e75da0_0 .net "temp_a_and_out", 0 0, L_0x5c7c3311d7d0;  1 drivers
v0x5c7c32e75f50_0 .net "temp_a_out", 0 0, L_0x5c7c3311d670;  1 drivers
v0x5c7c32e75ff0_0 .net "temp_b_and_out", 0 0, L_0x5c7c3311d9e0;  1 drivers
v0x5c7c32e761a0_0 .net "temp_b_out", 0 0, L_0x5c7c3311d880;  1 drivers
S_0x5c7c32e6bef0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e6bd10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e6cf90_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6d140_0 .net "in_b", 0 0, L_0x5c7c3311d670;  alias, 1 drivers
v0x5c7c32e6d230_0 .net "out", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
v0x5c7c32e6d350_0 .net "temp_out", 0 0, L_0x5c7c3311d720;  1 drivers
S_0x5c7c32e6c160 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e6bef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d720 .functor NAND 1, L_0x5c7c3311cfc0, L_0x5c7c3311d670, C4<1>, C4<1>;
v0x5c7c32e6c3d0_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6c490_0 .net "in_b", 0 0, L_0x5c7c3311d670;  alias, 1 drivers
v0x5c7c32e6c550_0 .net "out", 0 0, L_0x5c7c3311d720;  alias, 1 drivers
S_0x5c7c32e6c670 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e6bef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e6cde0_0 .net "in_a", 0 0, L_0x5c7c3311d720;  alias, 1 drivers
v0x5c7c32e6ce80_0 .net "out", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
S_0x5c7c32e6c890 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e6c670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d7d0 .functor NAND 1, L_0x5c7c3311d720, L_0x5c7c3311d720, C4<1>, C4<1>;
v0x5c7c32e6cb00_0 .net "in_a", 0 0, L_0x5c7c3311d720;  alias, 1 drivers
v0x5c7c32e6cbf0_0 .net "in_b", 0 0, L_0x5c7c3311d720;  alias, 1 drivers
v0x5c7c32e6cce0_0 .net "out", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
S_0x5c7c32e6d410 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e6bd10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e6e420_0 .net "in_a", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6e4c0_0 .net "in_b", 0 0, L_0x5c7c3311d880;  alias, 1 drivers
v0x5c7c32e6e5b0_0 .net "out", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
v0x5c7c32e6e6d0_0 .net "temp_out", 0 0, L_0x5c7c3311d930;  1 drivers
S_0x5c7c32e6d5f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e6d410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d930 .functor NAND 1, L_0x5c7c3311c0e0, L_0x5c7c3311d880, C4<1>, C4<1>;
v0x5c7c32e6d860_0 .net "in_a", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6d920_0 .net "in_b", 0 0, L_0x5c7c3311d880;  alias, 1 drivers
v0x5c7c32e6d9e0_0 .net "out", 0 0, L_0x5c7c3311d930;  alias, 1 drivers
S_0x5c7c32e6db00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e6d410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e6e270_0 .net "in_a", 0 0, L_0x5c7c3311d930;  alias, 1 drivers
v0x5c7c32e6e310_0 .net "out", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
S_0x5c7c32e6dd20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e6db00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d9e0 .functor NAND 1, L_0x5c7c3311d930, L_0x5c7c3311d930, C4<1>, C4<1>;
v0x5c7c32e6df90_0 .net "in_a", 0 0, L_0x5c7c3311d930;  alias, 1 drivers
v0x5c7c32e6e080_0 .net "in_b", 0 0, L_0x5c7c3311d930;  alias, 1 drivers
v0x5c7c32e6e170_0 .net "out", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
S_0x5c7c32e6e820 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e6bd10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e6f030_0 .net "in_a", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6f0d0_0 .net "out", 0 0, L_0x5c7c3311d670;  alias, 1 drivers
S_0x5c7c32e6e9f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e6e820;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d670 .functor NAND 1, L_0x5c7c3311c0e0, L_0x5c7c3311c0e0, C4<1>, C4<1>;
v0x5c7c32e6ec40_0 .net "in_a", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6ee10_0 .net "in_b", 0 0, L_0x5c7c3311c0e0;  alias, 1 drivers
v0x5c7c32e6eed0_0 .net "out", 0 0, L_0x5c7c3311d670;  alias, 1 drivers
S_0x5c7c32e6f1d0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e6bd10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e6f910_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6f9b0_0 .net "out", 0 0, L_0x5c7c3311d880;  alias, 1 drivers
S_0x5c7c32e6f3f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e6f1d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311d880 .functor NAND 1, L_0x5c7c3311cfc0, L_0x5c7c3311cfc0, C4<1>, C4<1>;
v0x5c7c32e6f660_0 .net "in_a", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6f720_0 .net "in_b", 0 0, L_0x5c7c3311cfc0;  alias, 1 drivers
v0x5c7c32e6f7e0_0 .net "out", 0 0, L_0x5c7c3311d880;  alias, 1 drivers
S_0x5c7c32e6fab0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e6bd10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e754f0_0 .net "branch1_out", 0 0, L_0x5c7c3311dbf0;  1 drivers
v0x5c7c32e75620_0 .net "branch2_out", 0 0, L_0x5c7c3311dd70;  1 drivers
v0x5c7c32e75770_0 .net "in_a", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
v0x5c7c32e75840_0 .net "in_b", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
v0x5c7c32e758e0_0 .net "out", 0 0, L_0x5c7c3311def0;  alias, 1 drivers
v0x5c7c32e75980_0 .net "temp1_out", 0 0, L_0x5c7c3311db40;  1 drivers
v0x5c7c32e75a20_0 .net "temp2_out", 0 0, L_0x5c7c3311dcc0;  1 drivers
v0x5c7c32e75ac0_0 .net "temp3_out", 0 0, L_0x5c7c3311de40;  1 drivers
S_0x5c7c32e6fd30 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e6fab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e70d30_0 .net "in_a", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
v0x5c7c32e70dd0_0 .net "in_b", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
v0x5c7c32e70e90_0 .net "out", 0 0, L_0x5c7c3311db40;  alias, 1 drivers
v0x5c7c32e70fb0_0 .net "temp_out", 0 0, L_0x5c7c3311da90;  1 drivers
S_0x5c7c32e6ffa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e6fd30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311da90 .functor NAND 1, L_0x5c7c3311d7d0, L_0x5c7c3311d7d0, C4<1>, C4<1>;
v0x5c7c32e70210_0 .net "in_a", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
v0x5c7c32e702d0_0 .net "in_b", 0 0, L_0x5c7c3311d7d0;  alias, 1 drivers
v0x5c7c32e70390_0 .net "out", 0 0, L_0x5c7c3311da90;  alias, 1 drivers
S_0x5c7c32e70490 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e6fd30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e70b80_0 .net "in_a", 0 0, L_0x5c7c3311da90;  alias, 1 drivers
v0x5c7c32e70c20_0 .net "out", 0 0, L_0x5c7c3311db40;  alias, 1 drivers
S_0x5c7c32e70660 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e70490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311db40 .functor NAND 1, L_0x5c7c3311da90, L_0x5c7c3311da90, C4<1>, C4<1>;
v0x5c7c32e708d0_0 .net "in_a", 0 0, L_0x5c7c3311da90;  alias, 1 drivers
v0x5c7c32e70990_0 .net "in_b", 0 0, L_0x5c7c3311da90;  alias, 1 drivers
v0x5c7c32e70a80_0 .net "out", 0 0, L_0x5c7c3311db40;  alias, 1 drivers
S_0x5c7c32e71120 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e6fab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e72150_0 .net "in_a", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
v0x5c7c32e721f0_0 .net "in_b", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
v0x5c7c32e722b0_0 .net "out", 0 0, L_0x5c7c3311dcc0;  alias, 1 drivers
v0x5c7c32e723d0_0 .net "temp_out", 0 0, L_0x5c7c32e73f70;  1 drivers
S_0x5c7c32e71300 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e71120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e73f70 .functor NAND 1, L_0x5c7c3311d9e0, L_0x5c7c3311d9e0, C4<1>, C4<1>;
v0x5c7c32e71570_0 .net "in_a", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
v0x5c7c32e71630_0 .net "in_b", 0 0, L_0x5c7c3311d9e0;  alias, 1 drivers
v0x5c7c32e71780_0 .net "out", 0 0, L_0x5c7c32e73f70;  alias, 1 drivers
S_0x5c7c32e71880 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e71120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e71fa0_0 .net "in_a", 0 0, L_0x5c7c32e73f70;  alias, 1 drivers
v0x5c7c32e72040_0 .net "out", 0 0, L_0x5c7c3311dcc0;  alias, 1 drivers
S_0x5c7c32e71a50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e71880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311dcc0 .functor NAND 1, L_0x5c7c32e73f70, L_0x5c7c32e73f70, C4<1>, C4<1>;
v0x5c7c32e71cc0_0 .net "in_a", 0 0, L_0x5c7c32e73f70;  alias, 1 drivers
v0x5c7c32e71db0_0 .net "in_b", 0 0, L_0x5c7c32e73f70;  alias, 1 drivers
v0x5c7c32e71ea0_0 .net "out", 0 0, L_0x5c7c3311dcc0;  alias, 1 drivers
S_0x5c7c32e72540 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e6fab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e73580_0 .net "in_a", 0 0, L_0x5c7c3311dbf0;  alias, 1 drivers
v0x5c7c32e73650_0 .net "in_b", 0 0, L_0x5c7c3311dd70;  alias, 1 drivers
v0x5c7c32e73720_0 .net "out", 0 0, L_0x5c7c3311de40;  alias, 1 drivers
v0x5c7c32e73840_0 .net "temp_out", 0 0, L_0x5c7c32e748e0;  1 drivers
S_0x5c7c32e72720 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e72540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e748e0 .functor NAND 1, L_0x5c7c3311dbf0, L_0x5c7c3311dd70, C4<1>, C4<1>;
v0x5c7c32e72970_0 .net "in_a", 0 0, L_0x5c7c3311dbf0;  alias, 1 drivers
v0x5c7c32e72a50_0 .net "in_b", 0 0, L_0x5c7c3311dd70;  alias, 1 drivers
v0x5c7c32e72b10_0 .net "out", 0 0, L_0x5c7c32e748e0;  alias, 1 drivers
S_0x5c7c32e72c60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e72540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e733d0_0 .net "in_a", 0 0, L_0x5c7c32e748e0;  alias, 1 drivers
v0x5c7c32e73470_0 .net "out", 0 0, L_0x5c7c3311de40;  alias, 1 drivers
S_0x5c7c32e72e80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e72c60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311de40 .functor NAND 1, L_0x5c7c32e748e0, L_0x5c7c32e748e0, C4<1>, C4<1>;
v0x5c7c32e730f0_0 .net "in_a", 0 0, L_0x5c7c32e748e0;  alias, 1 drivers
v0x5c7c32e731e0_0 .net "in_b", 0 0, L_0x5c7c32e748e0;  alias, 1 drivers
v0x5c7c32e732d0_0 .net "out", 0 0, L_0x5c7c3311de40;  alias, 1 drivers
S_0x5c7c32e73990 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e6fab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e740c0_0 .net "in_a", 0 0, L_0x5c7c3311db40;  alias, 1 drivers
v0x5c7c32e74160_0 .net "out", 0 0, L_0x5c7c3311dbf0;  alias, 1 drivers
S_0x5c7c32e73b60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e73990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311dbf0 .functor NAND 1, L_0x5c7c3311db40, L_0x5c7c3311db40, C4<1>, C4<1>;
v0x5c7c32e73dd0_0 .net "in_a", 0 0, L_0x5c7c3311db40;  alias, 1 drivers
v0x5c7c32e73e90_0 .net "in_b", 0 0, L_0x5c7c3311db40;  alias, 1 drivers
v0x5c7c32e73fe0_0 .net "out", 0 0, L_0x5c7c3311dbf0;  alias, 1 drivers
S_0x5c7c32e74260 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e6fab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e74a30_0 .net "in_a", 0 0, L_0x5c7c3311dcc0;  alias, 1 drivers
v0x5c7c32e74ad0_0 .net "out", 0 0, L_0x5c7c3311dd70;  alias, 1 drivers
S_0x5c7c32e744d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e74260;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311dd70 .functor NAND 1, L_0x5c7c3311dcc0, L_0x5c7c3311dcc0, C4<1>, C4<1>;
v0x5c7c32e74740_0 .net "in_a", 0 0, L_0x5c7c3311dcc0;  alias, 1 drivers
v0x5c7c32e74800_0 .net "in_b", 0 0, L_0x5c7c3311dcc0;  alias, 1 drivers
v0x5c7c32e74950_0 .net "out", 0 0, L_0x5c7c3311dd70;  alias, 1 drivers
S_0x5c7c32e74bd0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e6fab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e75370_0 .net "in_a", 0 0, L_0x5c7c3311de40;  alias, 1 drivers
v0x5c7c32e75410_0 .net "out", 0 0, L_0x5c7c3311def0;  alias, 1 drivers
S_0x5c7c32e74df0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e74bd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311def0 .functor NAND 1, L_0x5c7c3311de40, L_0x5c7c3311de40, C4<1>, C4<1>;
v0x5c7c32e75060_0 .net "in_a", 0 0, L_0x5c7c3311de40;  alias, 1 drivers
v0x5c7c32e75120_0 .net "in_b", 0 0, L_0x5c7c3311de40;  alias, 1 drivers
v0x5c7c32e75270_0 .net "out", 0 0, L_0x5c7c3311def0;  alias, 1 drivers
S_0x5c7c32e765f0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32e5e480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e7bfe0_0 .net "branch1_out", 0 0, L_0x5c7c3311e180;  1 drivers
v0x5c7c32e7c110_0 .net "branch2_out", 0 0, L_0x5c7c3311e410;  1 drivers
v0x5c7c32e7c260_0 .net "in_a", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e7c440_0 .net "in_b", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e7c5f0_0 .net "out", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e7c690_0 .net "temp1_out", 0 0, L_0x5c7c3311e0d0;  1 drivers
v0x5c7c32e7c730_0 .net "temp2_out", 0 0, L_0x5c7c3311e360;  1 drivers
v0x5c7c32e7c7d0_0 .net "temp3_out", 0 0, L_0x5c7c3311e5f0;  1 drivers
S_0x5c7c32e76780 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e765f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e77820_0 .net "in_a", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e778c0_0 .net "in_b", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e77980_0 .net "out", 0 0, L_0x5c7c3311e0d0;  alias, 1 drivers
v0x5c7c32e77aa0_0 .net "temp_out", 0 0, L_0x5c7c32e75200;  1 drivers
S_0x5c7c32e769a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e76780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e75200 .functor NAND 1, L_0x5c7c3311c470, L_0x5c7c3311c470, C4<1>, C4<1>;
v0x5c7c32e76c10_0 .net "in_a", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e76d60_0 .net "in_b", 0 0, L_0x5c7c3311c470;  alias, 1 drivers
v0x5c7c32e76e20_0 .net "out", 0 0, L_0x5c7c32e75200;  alias, 1 drivers
S_0x5c7c32e76f50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e76780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e77670_0 .net "in_a", 0 0, L_0x5c7c32e75200;  alias, 1 drivers
v0x5c7c32e77710_0 .net "out", 0 0, L_0x5c7c3311e0d0;  alias, 1 drivers
S_0x5c7c32e77120 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e76f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e0d0 .functor NAND 1, L_0x5c7c32e75200, L_0x5c7c32e75200, C4<1>, C4<1>;
v0x5c7c32e77390_0 .net "in_a", 0 0, L_0x5c7c32e75200;  alias, 1 drivers
v0x5c7c32e77480_0 .net "in_b", 0 0, L_0x5c7c32e75200;  alias, 1 drivers
v0x5c7c32e77570_0 .net "out", 0 0, L_0x5c7c3311e0d0;  alias, 1 drivers
S_0x5c7c32e77c10 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e765f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e78c40_0 .net "in_a", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e78ce0_0 .net "in_b", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e78da0_0 .net "out", 0 0, L_0x5c7c3311e360;  alias, 1 drivers
v0x5c7c32e78ec0_0 .net "temp_out", 0 0, L_0x5c7c32e7aa60;  1 drivers
S_0x5c7c32e77df0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e77c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e7aa60 .functor NAND 1, L_0x5c7c3311d5c0, L_0x5c7c3311d5c0, C4<1>, C4<1>;
v0x5c7c32e78060_0 .net "in_a", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e781b0_0 .net "in_b", 0 0, L_0x5c7c3311d5c0;  alias, 1 drivers
v0x5c7c32e78270_0 .net "out", 0 0, L_0x5c7c32e7aa60;  alias, 1 drivers
S_0x5c7c32e78370 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e77c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e78a90_0 .net "in_a", 0 0, L_0x5c7c32e7aa60;  alias, 1 drivers
v0x5c7c32e78b30_0 .net "out", 0 0, L_0x5c7c3311e360;  alias, 1 drivers
S_0x5c7c32e78540 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e78370;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e360 .functor NAND 1, L_0x5c7c32e7aa60, L_0x5c7c32e7aa60, C4<1>, C4<1>;
v0x5c7c32e787b0_0 .net "in_a", 0 0, L_0x5c7c32e7aa60;  alias, 1 drivers
v0x5c7c32e788a0_0 .net "in_b", 0 0, L_0x5c7c32e7aa60;  alias, 1 drivers
v0x5c7c32e78990_0 .net "out", 0 0, L_0x5c7c3311e360;  alias, 1 drivers
S_0x5c7c32e79030 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e765f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e7a070_0 .net "in_a", 0 0, L_0x5c7c3311e180;  alias, 1 drivers
v0x5c7c32e7a140_0 .net "in_b", 0 0, L_0x5c7c3311e410;  alias, 1 drivers
v0x5c7c32e7a210_0 .net "out", 0 0, L_0x5c7c3311e5f0;  alias, 1 drivers
v0x5c7c32e7a330_0 .net "temp_out", 0 0, L_0x5c7c32e7b3d0;  1 drivers
S_0x5c7c32e79210 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e79030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e7b3d0 .functor NAND 1, L_0x5c7c3311e180, L_0x5c7c3311e410, C4<1>, C4<1>;
v0x5c7c32e79460_0 .net "in_a", 0 0, L_0x5c7c3311e180;  alias, 1 drivers
v0x5c7c32e79540_0 .net "in_b", 0 0, L_0x5c7c3311e410;  alias, 1 drivers
v0x5c7c32e79600_0 .net "out", 0 0, L_0x5c7c32e7b3d0;  alias, 1 drivers
S_0x5c7c32e79750 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e79030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e79ec0_0 .net "in_a", 0 0, L_0x5c7c32e7b3d0;  alias, 1 drivers
v0x5c7c32e79f60_0 .net "out", 0 0, L_0x5c7c3311e5f0;  alias, 1 drivers
S_0x5c7c32e79970 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e79750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e5f0 .functor NAND 1, L_0x5c7c32e7b3d0, L_0x5c7c32e7b3d0, C4<1>, C4<1>;
v0x5c7c32e79be0_0 .net "in_a", 0 0, L_0x5c7c32e7b3d0;  alias, 1 drivers
v0x5c7c32e79cd0_0 .net "in_b", 0 0, L_0x5c7c32e7b3d0;  alias, 1 drivers
v0x5c7c32e79dc0_0 .net "out", 0 0, L_0x5c7c3311e5f0;  alias, 1 drivers
S_0x5c7c32e7a480 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e765f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e7abb0_0 .net "in_a", 0 0, L_0x5c7c3311e0d0;  alias, 1 drivers
v0x5c7c32e7ac50_0 .net "out", 0 0, L_0x5c7c3311e180;  alias, 1 drivers
S_0x5c7c32e7a650 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e7a480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e180 .functor NAND 1, L_0x5c7c3311e0d0, L_0x5c7c3311e0d0, C4<1>, C4<1>;
v0x5c7c32e7a8c0_0 .net "in_a", 0 0, L_0x5c7c3311e0d0;  alias, 1 drivers
v0x5c7c32e7a980_0 .net "in_b", 0 0, L_0x5c7c3311e0d0;  alias, 1 drivers
v0x5c7c32e7aad0_0 .net "out", 0 0, L_0x5c7c3311e180;  alias, 1 drivers
S_0x5c7c32e7ad50 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e765f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e7b520_0 .net "in_a", 0 0, L_0x5c7c3311e360;  alias, 1 drivers
v0x5c7c32e7b5c0_0 .net "out", 0 0, L_0x5c7c3311e410;  alias, 1 drivers
S_0x5c7c32e7afc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e7ad50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e410 .functor NAND 1, L_0x5c7c3311e360, L_0x5c7c3311e360, C4<1>, C4<1>;
v0x5c7c32e7b230_0 .net "in_a", 0 0, L_0x5c7c3311e360;  alias, 1 drivers
v0x5c7c32e7b2f0_0 .net "in_b", 0 0, L_0x5c7c3311e360;  alias, 1 drivers
v0x5c7c32e7b440_0 .net "out", 0 0, L_0x5c7c3311e410;  alias, 1 drivers
S_0x5c7c32e7b6c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e765f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e7be60_0 .net "in_a", 0 0, L_0x5c7c3311e5f0;  alias, 1 drivers
v0x5c7c32e7bf00_0 .net "out", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
S_0x5c7c32e7b8e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e7b6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e6a0 .functor NAND 1, L_0x5c7c3311e5f0, L_0x5c7c3311e5f0, C4<1>, C4<1>;
v0x5c7c32e7bb50_0 .net "in_a", 0 0, L_0x5c7c3311e5f0;  alias, 1 drivers
v0x5c7c32e7bc10_0 .net "in_b", 0 0, L_0x5c7c3311e5f0;  alias, 1 drivers
v0x5c7c32e7bd60_0 .net "out", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
S_0x5c7c32e7ce30 .scope module, "fa_gate7" "FullAdder" 2 12, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32e9b260_0 .net "a", 0 0, L_0x5c7c33120d90;  1 drivers
v0x5c7c32e9b300_0 .net "b", 0 0, L_0x5c7c33120e30;  1 drivers
v0x5c7c32e9b3c0_0 .net "c", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e9b460_0 .net "carry", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32e9b500_0 .net "sum", 0 0, L_0x5c7c33120440;  1 drivers
v0x5c7c32e9b5a0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c3311e9c0;  1 drivers
v0x5c7c32e9b640_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c3311fb10;  1 drivers
v0x5c7c32e9b6e0_0 .net "tmp_sum_out", 0 0, L_0x5c7c3311f510;  1 drivers
S_0x5c7c32e7d090 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32e7ce30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e88c10_0 .net "a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e88dc0_0 .net "b", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e88f90_0 .net "carry", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e89030_0 .net "sum", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
S_0x5c7c32e7d300 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e7d090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e7e3f0_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e7e4c0_0 .net "in_b", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e7e590_0 .net "out", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e7e6b0_0 .net "temp_out", 0 0, L_0x5c7c32e7bcf0;  1 drivers
S_0x5c7c32e7d570 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e7d300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e7bcf0 .functor NAND 1, L_0x5c7c33120d90, L_0x5c7c33120e30, C4<1>, C4<1>;
v0x5c7c32e7d7e0_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e7d8c0_0 .net "in_b", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e7d980_0 .net "out", 0 0, L_0x5c7c32e7bcf0;  alias, 1 drivers
S_0x5c7c32e7dad0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e7d300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e7e240_0 .net "in_a", 0 0, L_0x5c7c32e7bcf0;  alias, 1 drivers
v0x5c7c32e7e2e0_0 .net "out", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
S_0x5c7c32e7dcf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e7dad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311e9c0 .functor NAND 1, L_0x5c7c32e7bcf0, L_0x5c7c32e7bcf0, C4<1>, C4<1>;
v0x5c7c32e7df60_0 .net "in_a", 0 0, L_0x5c7c32e7bcf0;  alias, 1 drivers
v0x5c7c32e7e050_0 .net "in_b", 0 0, L_0x5c7c32e7bcf0;  alias, 1 drivers
v0x5c7c32e7e140_0 .net "out", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
S_0x5c7c32e7e770 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e7d090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e88530_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e885d0_0 .net "in_b", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e88690_0 .net "out", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e88730_0 .net "temp_a_and_out", 0 0, L_0x5c7c3311ebd0;  1 drivers
v0x5c7c32e888e0_0 .net "temp_a_out", 0 0, L_0x5c7c3311ea70;  1 drivers
v0x5c7c32e88980_0 .net "temp_b_and_out", 0 0, L_0x5c7c3311ede0;  1 drivers
v0x5c7c32e88b30_0 .net "temp_b_out", 0 0, L_0x5c7c3311ec80;  1 drivers
S_0x5c7c32e7e950 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e7e770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e7fa10_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e7fab0_0 .net "in_b", 0 0, L_0x5c7c3311ea70;  alias, 1 drivers
v0x5c7c32e7fba0_0 .net "out", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
v0x5c7c32e7fcc0_0 .net "temp_out", 0 0, L_0x5c7c3311eb20;  1 drivers
S_0x5c7c32e7ebc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e7e950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311eb20 .functor NAND 1, L_0x5c7c33120d90, L_0x5c7c3311ea70, C4<1>, C4<1>;
v0x5c7c32e7ee30_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e7ef40_0 .net "in_b", 0 0, L_0x5c7c3311ea70;  alias, 1 drivers
v0x5c7c32e7f000_0 .net "out", 0 0, L_0x5c7c3311eb20;  alias, 1 drivers
S_0x5c7c32e7f120 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e7e950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e7f860_0 .net "in_a", 0 0, L_0x5c7c3311eb20;  alias, 1 drivers
v0x5c7c32e7f900_0 .net "out", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
S_0x5c7c32e7f340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e7f120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ebd0 .functor NAND 1, L_0x5c7c3311eb20, L_0x5c7c3311eb20, C4<1>, C4<1>;
v0x5c7c32e7f5b0_0 .net "in_a", 0 0, L_0x5c7c3311eb20;  alias, 1 drivers
v0x5c7c32e7f670_0 .net "in_b", 0 0, L_0x5c7c3311eb20;  alias, 1 drivers
v0x5c7c32e7f760_0 .net "out", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
S_0x5c7c32e7fd80 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e7e770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e80db0_0 .net "in_a", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e80e50_0 .net "in_b", 0 0, L_0x5c7c3311ec80;  alias, 1 drivers
v0x5c7c32e80f40_0 .net "out", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
v0x5c7c32e81060_0 .net "temp_out", 0 0, L_0x5c7c3311ed30;  1 drivers
S_0x5c7c32e7ff60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e7fd80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ed30 .functor NAND 1, L_0x5c7c33120e30, L_0x5c7c3311ec80, C4<1>, C4<1>;
v0x5c7c32e801d0_0 .net "in_a", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e802e0_0 .net "in_b", 0 0, L_0x5c7c3311ec80;  alias, 1 drivers
v0x5c7c32e803a0_0 .net "out", 0 0, L_0x5c7c3311ed30;  alias, 1 drivers
S_0x5c7c32e804c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e7fd80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e80c00_0 .net "in_a", 0 0, L_0x5c7c3311ed30;  alias, 1 drivers
v0x5c7c32e80ca0_0 .net "out", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
S_0x5c7c32e806e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e804c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ede0 .functor NAND 1, L_0x5c7c3311ed30, L_0x5c7c3311ed30, C4<1>, C4<1>;
v0x5c7c32e80950_0 .net "in_a", 0 0, L_0x5c7c3311ed30;  alias, 1 drivers
v0x5c7c32e80a10_0 .net "in_b", 0 0, L_0x5c7c3311ed30;  alias, 1 drivers
v0x5c7c32e80b00_0 .net "out", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
S_0x5c7c32e811b0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e7e770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e818f0_0 .net "in_a", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e81990_0 .net "out", 0 0, L_0x5c7c3311ea70;  alias, 1 drivers
S_0x5c7c32e81380 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e811b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ea70 .functor NAND 1, L_0x5c7c33120e30, L_0x5c7c33120e30, C4<1>, C4<1>;
v0x5c7c32e815d0_0 .net "in_a", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e81720_0 .net "in_b", 0 0, L_0x5c7c33120e30;  alias, 1 drivers
v0x5c7c32e817e0_0 .net "out", 0 0, L_0x5c7c3311ea70;  alias, 1 drivers
S_0x5c7c32e81a90 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e7e770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e82210_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e822b0_0 .net "out", 0 0, L_0x5c7c3311ec80;  alias, 1 drivers
S_0x5c7c32e81cb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e81a90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ec80 .functor NAND 1, L_0x5c7c33120d90, L_0x5c7c33120d90, C4<1>, C4<1>;
v0x5c7c32e81f20_0 .net "in_a", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e82070_0 .net "in_b", 0 0, L_0x5c7c33120d90;  alias, 1 drivers
v0x5c7c32e82130_0 .net "out", 0 0, L_0x5c7c3311ec80;  alias, 1 drivers
S_0x5c7c32e823b0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e7e770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e87e80_0 .net "branch1_out", 0 0, L_0x5c7c3311eff0;  1 drivers
v0x5c7c32e87fb0_0 .net "branch2_out", 0 0, L_0x5c7c3311f280;  1 drivers
v0x5c7c32e88100_0 .net "in_a", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
v0x5c7c32e881d0_0 .net "in_b", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
v0x5c7c32e88270_0 .net "out", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e88310_0 .net "temp1_out", 0 0, L_0x5c7c3311ef40;  1 drivers
v0x5c7c32e883b0_0 .net "temp2_out", 0 0, L_0x5c7c3311f1d0;  1 drivers
v0x5c7c32e88450_0 .net "temp3_out", 0 0, L_0x5c7c3311f460;  1 drivers
S_0x5c7c32e82630 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e823b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e836c0_0 .net "in_a", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
v0x5c7c32e83760_0 .net "in_b", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
v0x5c7c32e83820_0 .net "out", 0 0, L_0x5c7c3311ef40;  alias, 1 drivers
v0x5c7c32e83940_0 .net "temp_out", 0 0, L_0x5c7c3311ee90;  1 drivers
S_0x5c7c32e828a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e82630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ee90 .functor NAND 1, L_0x5c7c3311ebd0, L_0x5c7c3311ebd0, C4<1>, C4<1>;
v0x5c7c32e82b10_0 .net "in_a", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
v0x5c7c32e82bd0_0 .net "in_b", 0 0, L_0x5c7c3311ebd0;  alias, 1 drivers
v0x5c7c32e82d20_0 .net "out", 0 0, L_0x5c7c3311ee90;  alias, 1 drivers
S_0x5c7c32e82e20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e82630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e83510_0 .net "in_a", 0 0, L_0x5c7c3311ee90;  alias, 1 drivers
v0x5c7c32e835b0_0 .net "out", 0 0, L_0x5c7c3311ef40;  alias, 1 drivers
S_0x5c7c32e82ff0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e82e20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ef40 .functor NAND 1, L_0x5c7c3311ee90, L_0x5c7c3311ee90, C4<1>, C4<1>;
v0x5c7c32e83260_0 .net "in_a", 0 0, L_0x5c7c3311ee90;  alias, 1 drivers
v0x5c7c32e83320_0 .net "in_b", 0 0, L_0x5c7c3311ee90;  alias, 1 drivers
v0x5c7c32e83410_0 .net "out", 0 0, L_0x5c7c3311ef40;  alias, 1 drivers
S_0x5c7c32e83ab0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e823b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e84ae0_0 .net "in_a", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
v0x5c7c32e84b80_0 .net "in_b", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
v0x5c7c32e84c40_0 .net "out", 0 0, L_0x5c7c3311f1d0;  alias, 1 drivers
v0x5c7c32e84d60_0 .net "temp_out", 0 0, L_0x5c7c32e86900;  1 drivers
S_0x5c7c32e83c90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e83ab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e86900 .functor NAND 1, L_0x5c7c3311ede0, L_0x5c7c3311ede0, C4<1>, C4<1>;
v0x5c7c32e83f00_0 .net "in_a", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
v0x5c7c32e83fc0_0 .net "in_b", 0 0, L_0x5c7c3311ede0;  alias, 1 drivers
v0x5c7c32e84110_0 .net "out", 0 0, L_0x5c7c32e86900;  alias, 1 drivers
S_0x5c7c32e84210 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e83ab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e84930_0 .net "in_a", 0 0, L_0x5c7c32e86900;  alias, 1 drivers
v0x5c7c32e849d0_0 .net "out", 0 0, L_0x5c7c3311f1d0;  alias, 1 drivers
S_0x5c7c32e843e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e84210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311f1d0 .functor NAND 1, L_0x5c7c32e86900, L_0x5c7c32e86900, C4<1>, C4<1>;
v0x5c7c32e84650_0 .net "in_a", 0 0, L_0x5c7c32e86900;  alias, 1 drivers
v0x5c7c32e84740_0 .net "in_b", 0 0, L_0x5c7c32e86900;  alias, 1 drivers
v0x5c7c32e84830_0 .net "out", 0 0, L_0x5c7c3311f1d0;  alias, 1 drivers
S_0x5c7c32e84ed0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e823b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e85f10_0 .net "in_a", 0 0, L_0x5c7c3311eff0;  alias, 1 drivers
v0x5c7c32e85fe0_0 .net "in_b", 0 0, L_0x5c7c3311f280;  alias, 1 drivers
v0x5c7c32e860b0_0 .net "out", 0 0, L_0x5c7c3311f460;  alias, 1 drivers
v0x5c7c32e861d0_0 .net "temp_out", 0 0, L_0x5c7c32e87270;  1 drivers
S_0x5c7c32e850b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e84ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e87270 .functor NAND 1, L_0x5c7c3311eff0, L_0x5c7c3311f280, C4<1>, C4<1>;
v0x5c7c32e85300_0 .net "in_a", 0 0, L_0x5c7c3311eff0;  alias, 1 drivers
v0x5c7c32e853e0_0 .net "in_b", 0 0, L_0x5c7c3311f280;  alias, 1 drivers
v0x5c7c32e854a0_0 .net "out", 0 0, L_0x5c7c32e87270;  alias, 1 drivers
S_0x5c7c32e855f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e84ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e85d60_0 .net "in_a", 0 0, L_0x5c7c32e87270;  alias, 1 drivers
v0x5c7c32e85e00_0 .net "out", 0 0, L_0x5c7c3311f460;  alias, 1 drivers
S_0x5c7c32e85810 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e855f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311f460 .functor NAND 1, L_0x5c7c32e87270, L_0x5c7c32e87270, C4<1>, C4<1>;
v0x5c7c32e85a80_0 .net "in_a", 0 0, L_0x5c7c32e87270;  alias, 1 drivers
v0x5c7c32e85b70_0 .net "in_b", 0 0, L_0x5c7c32e87270;  alias, 1 drivers
v0x5c7c32e85c60_0 .net "out", 0 0, L_0x5c7c3311f460;  alias, 1 drivers
S_0x5c7c32e86320 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e823b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e86a50_0 .net "in_a", 0 0, L_0x5c7c3311ef40;  alias, 1 drivers
v0x5c7c32e86af0_0 .net "out", 0 0, L_0x5c7c3311eff0;  alias, 1 drivers
S_0x5c7c32e864f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e86320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311eff0 .functor NAND 1, L_0x5c7c3311ef40, L_0x5c7c3311ef40, C4<1>, C4<1>;
v0x5c7c32e86760_0 .net "in_a", 0 0, L_0x5c7c3311ef40;  alias, 1 drivers
v0x5c7c32e86820_0 .net "in_b", 0 0, L_0x5c7c3311ef40;  alias, 1 drivers
v0x5c7c32e86970_0 .net "out", 0 0, L_0x5c7c3311eff0;  alias, 1 drivers
S_0x5c7c32e86bf0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e823b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e873c0_0 .net "in_a", 0 0, L_0x5c7c3311f1d0;  alias, 1 drivers
v0x5c7c32e87460_0 .net "out", 0 0, L_0x5c7c3311f280;  alias, 1 drivers
S_0x5c7c32e86e60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e86bf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311f280 .functor NAND 1, L_0x5c7c3311f1d0, L_0x5c7c3311f1d0, C4<1>, C4<1>;
v0x5c7c32e870d0_0 .net "in_a", 0 0, L_0x5c7c3311f1d0;  alias, 1 drivers
v0x5c7c32e87190_0 .net "in_b", 0 0, L_0x5c7c3311f1d0;  alias, 1 drivers
v0x5c7c32e872e0_0 .net "out", 0 0, L_0x5c7c3311f280;  alias, 1 drivers
S_0x5c7c32e87560 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e823b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e87d00_0 .net "in_a", 0 0, L_0x5c7c3311f460;  alias, 1 drivers
v0x5c7c32e87da0_0 .net "out", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
S_0x5c7c32e87780 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e87560;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311f510 .functor NAND 1, L_0x5c7c3311f460, L_0x5c7c3311f460, C4<1>, C4<1>;
v0x5c7c32e879f0_0 .net "in_a", 0 0, L_0x5c7c3311f460;  alias, 1 drivers
v0x5c7c32e87ab0_0 .net "in_b", 0 0, L_0x5c7c3311f460;  alias, 1 drivers
v0x5c7c32e87c00_0 .net "out", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
S_0x5c7c32e89110 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32e7ce30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32e94c30_0 .net "a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e94cd0_0 .net "b", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e94d90_0 .net "carry", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e94e30_0 .net "sum", 0 0, L_0x5c7c33120440;  alias, 1 drivers
S_0x5c7c32e89330 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e89110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e8a2d0_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e8a370_0 .net "in_b", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e8a430_0 .net "out", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e8a550_0 .net "temp_out", 0 0, L_0x5c7c32e87b90;  1 drivers
S_0x5c7c32e894e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e89330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e87b90 .functor NAND 1, L_0x5c7c3311f510, L_0x5c7c3311e6a0, C4<1>, C4<1>;
v0x5c7c32e89750_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e89810_0 .net "in_b", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e898d0_0 .net "out", 0 0, L_0x5c7c32e87b90;  alias, 1 drivers
S_0x5c7c32e89a00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e89330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e8a120_0 .net "in_a", 0 0, L_0x5c7c32e87b90;  alias, 1 drivers
v0x5c7c32e8a1c0_0 .net "out", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
S_0x5c7c32e89bd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e89a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311fb10 .functor NAND 1, L_0x5c7c32e87b90, L_0x5c7c32e87b90, C4<1>, C4<1>;
v0x5c7c32e89e40_0 .net "in_a", 0 0, L_0x5c7c32e87b90;  alias, 1 drivers
v0x5c7c32e89f30_0 .net "in_b", 0 0, L_0x5c7c32e87b90;  alias, 1 drivers
v0x5c7c32e8a020_0 .net "out", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
S_0x5c7c32e8a6c0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e89110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e94550_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e945f0_0 .net "in_b", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e946b0_0 .net "out", 0 0, L_0x5c7c33120440;  alias, 1 drivers
v0x5c7c32e94750_0 .net "temp_a_and_out", 0 0, L_0x5c7c3311fd20;  1 drivers
v0x5c7c32e94900_0 .net "temp_a_out", 0 0, L_0x5c7c3311fbc0;  1 drivers
v0x5c7c32e949a0_0 .net "temp_b_and_out", 0 0, L_0x5c7c3311ff30;  1 drivers
v0x5c7c32e94b50_0 .net "temp_b_out", 0 0, L_0x5c7c3311fdd0;  1 drivers
S_0x5c7c32e8a8a0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e8a6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e8b940_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e8baf0_0 .net "in_b", 0 0, L_0x5c7c3311fbc0;  alias, 1 drivers
v0x5c7c32e8bbe0_0 .net "out", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
v0x5c7c32e8bd00_0 .net "temp_out", 0 0, L_0x5c7c3311fc70;  1 drivers
S_0x5c7c32e8ab10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e8a8a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311fc70 .functor NAND 1, L_0x5c7c3311f510, L_0x5c7c3311fbc0, C4<1>, C4<1>;
v0x5c7c32e8ad80_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e8ae40_0 .net "in_b", 0 0, L_0x5c7c3311fbc0;  alias, 1 drivers
v0x5c7c32e8af00_0 .net "out", 0 0, L_0x5c7c3311fc70;  alias, 1 drivers
S_0x5c7c32e8b020 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e8a8a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e8b790_0 .net "in_a", 0 0, L_0x5c7c3311fc70;  alias, 1 drivers
v0x5c7c32e8b830_0 .net "out", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
S_0x5c7c32e8b240 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e8b020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311fd20 .functor NAND 1, L_0x5c7c3311fc70, L_0x5c7c3311fc70, C4<1>, C4<1>;
v0x5c7c32e8b4b0_0 .net "in_a", 0 0, L_0x5c7c3311fc70;  alias, 1 drivers
v0x5c7c32e8b5a0_0 .net "in_b", 0 0, L_0x5c7c3311fc70;  alias, 1 drivers
v0x5c7c32e8b690_0 .net "out", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
S_0x5c7c32e8bdc0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e8a6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e8cdd0_0 .net "in_a", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e8ce70_0 .net "in_b", 0 0, L_0x5c7c3311fdd0;  alias, 1 drivers
v0x5c7c32e8cf60_0 .net "out", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
v0x5c7c32e8d080_0 .net "temp_out", 0 0, L_0x5c7c3311fe80;  1 drivers
S_0x5c7c32e8bfa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e8bdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311fe80 .functor NAND 1, L_0x5c7c3311e6a0, L_0x5c7c3311fdd0, C4<1>, C4<1>;
v0x5c7c32e8c210_0 .net "in_a", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e8c2d0_0 .net "in_b", 0 0, L_0x5c7c3311fdd0;  alias, 1 drivers
v0x5c7c32e8c390_0 .net "out", 0 0, L_0x5c7c3311fe80;  alias, 1 drivers
S_0x5c7c32e8c4b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e8bdc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e8cc20_0 .net "in_a", 0 0, L_0x5c7c3311fe80;  alias, 1 drivers
v0x5c7c32e8ccc0_0 .net "out", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
S_0x5c7c32e8c6d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e8c4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ff30 .functor NAND 1, L_0x5c7c3311fe80, L_0x5c7c3311fe80, C4<1>, C4<1>;
v0x5c7c32e8c940_0 .net "in_a", 0 0, L_0x5c7c3311fe80;  alias, 1 drivers
v0x5c7c32e8ca30_0 .net "in_b", 0 0, L_0x5c7c3311fe80;  alias, 1 drivers
v0x5c7c32e8cb20_0 .net "out", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
S_0x5c7c32e8d1d0 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e8a6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e8d9e0_0 .net "in_a", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e8da80_0 .net "out", 0 0, L_0x5c7c3311fbc0;  alias, 1 drivers
S_0x5c7c32e8d3a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e8d1d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311fbc0 .functor NAND 1, L_0x5c7c3311e6a0, L_0x5c7c3311e6a0, C4<1>, C4<1>;
v0x5c7c32e8d5f0_0 .net "in_a", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e8d7c0_0 .net "in_b", 0 0, L_0x5c7c3311e6a0;  alias, 1 drivers
v0x5c7c32e8d880_0 .net "out", 0 0, L_0x5c7c3311fbc0;  alias, 1 drivers
S_0x5c7c32e8db80 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e8a6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e8e2c0_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e8e360_0 .net "out", 0 0, L_0x5c7c3311fdd0;  alias, 1 drivers
S_0x5c7c32e8dda0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e8db80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311fdd0 .functor NAND 1, L_0x5c7c3311f510, L_0x5c7c3311f510, C4<1>, C4<1>;
v0x5c7c32e8e010_0 .net "in_a", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e8e0d0_0 .net "in_b", 0 0, L_0x5c7c3311f510;  alias, 1 drivers
v0x5c7c32e8e190_0 .net "out", 0 0, L_0x5c7c3311fdd0;  alias, 1 drivers
S_0x5c7c32e8e460 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e8a6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e93ea0_0 .net "branch1_out", 0 0, L_0x5c7c33120140;  1 drivers
v0x5c7c32e93fd0_0 .net "branch2_out", 0 0, L_0x5c7c331202c0;  1 drivers
v0x5c7c32e94120_0 .net "in_a", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
v0x5c7c32e941f0_0 .net "in_b", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
v0x5c7c32e94290_0 .net "out", 0 0, L_0x5c7c33120440;  alias, 1 drivers
v0x5c7c32e94330_0 .net "temp1_out", 0 0, L_0x5c7c33120090;  1 drivers
v0x5c7c32e943d0_0 .net "temp2_out", 0 0, L_0x5c7c33120210;  1 drivers
v0x5c7c32e94470_0 .net "temp3_out", 0 0, L_0x5c7c33120390;  1 drivers
S_0x5c7c32e8e6e0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e8e460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e8f6e0_0 .net "in_a", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
v0x5c7c32e8f780_0 .net "in_b", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
v0x5c7c32e8f840_0 .net "out", 0 0, L_0x5c7c33120090;  alias, 1 drivers
v0x5c7c32e8f960_0 .net "temp_out", 0 0, L_0x5c7c3311ffe0;  1 drivers
S_0x5c7c32e8e950 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e8e6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3311ffe0 .functor NAND 1, L_0x5c7c3311fd20, L_0x5c7c3311fd20, C4<1>, C4<1>;
v0x5c7c32e8ebc0_0 .net "in_a", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
v0x5c7c32e8ec80_0 .net "in_b", 0 0, L_0x5c7c3311fd20;  alias, 1 drivers
v0x5c7c32e8ed40_0 .net "out", 0 0, L_0x5c7c3311ffe0;  alias, 1 drivers
S_0x5c7c32e8ee40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e8e6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e8f530_0 .net "in_a", 0 0, L_0x5c7c3311ffe0;  alias, 1 drivers
v0x5c7c32e8f5d0_0 .net "out", 0 0, L_0x5c7c33120090;  alias, 1 drivers
S_0x5c7c32e8f010 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e8ee40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120090 .functor NAND 1, L_0x5c7c3311ffe0, L_0x5c7c3311ffe0, C4<1>, C4<1>;
v0x5c7c32e8f280_0 .net "in_a", 0 0, L_0x5c7c3311ffe0;  alias, 1 drivers
v0x5c7c32e8f340_0 .net "in_b", 0 0, L_0x5c7c3311ffe0;  alias, 1 drivers
v0x5c7c32e8f430_0 .net "out", 0 0, L_0x5c7c33120090;  alias, 1 drivers
S_0x5c7c32e8fad0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e8e460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e90b00_0 .net "in_a", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
v0x5c7c32e90ba0_0 .net "in_b", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
v0x5c7c32e90c60_0 .net "out", 0 0, L_0x5c7c33120210;  alias, 1 drivers
v0x5c7c32e90d80_0 .net "temp_out", 0 0, L_0x5c7c32e92920;  1 drivers
S_0x5c7c32e8fcb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e8fad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e92920 .functor NAND 1, L_0x5c7c3311ff30, L_0x5c7c3311ff30, C4<1>, C4<1>;
v0x5c7c32e8ff20_0 .net "in_a", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
v0x5c7c32e8ffe0_0 .net "in_b", 0 0, L_0x5c7c3311ff30;  alias, 1 drivers
v0x5c7c32e90130_0 .net "out", 0 0, L_0x5c7c32e92920;  alias, 1 drivers
S_0x5c7c32e90230 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e8fad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e90950_0 .net "in_a", 0 0, L_0x5c7c32e92920;  alias, 1 drivers
v0x5c7c32e909f0_0 .net "out", 0 0, L_0x5c7c33120210;  alias, 1 drivers
S_0x5c7c32e90400 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e90230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120210 .functor NAND 1, L_0x5c7c32e92920, L_0x5c7c32e92920, C4<1>, C4<1>;
v0x5c7c32e90670_0 .net "in_a", 0 0, L_0x5c7c32e92920;  alias, 1 drivers
v0x5c7c32e90760_0 .net "in_b", 0 0, L_0x5c7c32e92920;  alias, 1 drivers
v0x5c7c32e90850_0 .net "out", 0 0, L_0x5c7c33120210;  alias, 1 drivers
S_0x5c7c32e90ef0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e8e460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e91f30_0 .net "in_a", 0 0, L_0x5c7c33120140;  alias, 1 drivers
v0x5c7c32e92000_0 .net "in_b", 0 0, L_0x5c7c331202c0;  alias, 1 drivers
v0x5c7c32e920d0_0 .net "out", 0 0, L_0x5c7c33120390;  alias, 1 drivers
v0x5c7c32e921f0_0 .net "temp_out", 0 0, L_0x5c7c32e93290;  1 drivers
S_0x5c7c32e910d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e90ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e93290 .functor NAND 1, L_0x5c7c33120140, L_0x5c7c331202c0, C4<1>, C4<1>;
v0x5c7c32e91320_0 .net "in_a", 0 0, L_0x5c7c33120140;  alias, 1 drivers
v0x5c7c32e91400_0 .net "in_b", 0 0, L_0x5c7c331202c0;  alias, 1 drivers
v0x5c7c32e914c0_0 .net "out", 0 0, L_0x5c7c32e93290;  alias, 1 drivers
S_0x5c7c32e91610 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e90ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e91d80_0 .net "in_a", 0 0, L_0x5c7c32e93290;  alias, 1 drivers
v0x5c7c32e91e20_0 .net "out", 0 0, L_0x5c7c33120390;  alias, 1 drivers
S_0x5c7c32e91830 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e91610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120390 .functor NAND 1, L_0x5c7c32e93290, L_0x5c7c32e93290, C4<1>, C4<1>;
v0x5c7c32e91aa0_0 .net "in_a", 0 0, L_0x5c7c32e93290;  alias, 1 drivers
v0x5c7c32e91b90_0 .net "in_b", 0 0, L_0x5c7c32e93290;  alias, 1 drivers
v0x5c7c32e91c80_0 .net "out", 0 0, L_0x5c7c33120390;  alias, 1 drivers
S_0x5c7c32e92340 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e8e460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e92a70_0 .net "in_a", 0 0, L_0x5c7c33120090;  alias, 1 drivers
v0x5c7c32e92b10_0 .net "out", 0 0, L_0x5c7c33120140;  alias, 1 drivers
S_0x5c7c32e92510 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e92340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120140 .functor NAND 1, L_0x5c7c33120090, L_0x5c7c33120090, C4<1>, C4<1>;
v0x5c7c32e92780_0 .net "in_a", 0 0, L_0x5c7c33120090;  alias, 1 drivers
v0x5c7c32e92840_0 .net "in_b", 0 0, L_0x5c7c33120090;  alias, 1 drivers
v0x5c7c32e92990_0 .net "out", 0 0, L_0x5c7c33120140;  alias, 1 drivers
S_0x5c7c32e92c10 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e8e460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e933e0_0 .net "in_a", 0 0, L_0x5c7c33120210;  alias, 1 drivers
v0x5c7c32e93480_0 .net "out", 0 0, L_0x5c7c331202c0;  alias, 1 drivers
S_0x5c7c32e92e80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e92c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331202c0 .functor NAND 1, L_0x5c7c33120210, L_0x5c7c33120210, C4<1>, C4<1>;
v0x5c7c32e930f0_0 .net "in_a", 0 0, L_0x5c7c33120210;  alias, 1 drivers
v0x5c7c32e931b0_0 .net "in_b", 0 0, L_0x5c7c33120210;  alias, 1 drivers
v0x5c7c32e93300_0 .net "out", 0 0, L_0x5c7c331202c0;  alias, 1 drivers
S_0x5c7c32e93580 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e8e460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e93d20_0 .net "in_a", 0 0, L_0x5c7c33120390;  alias, 1 drivers
v0x5c7c32e93dc0_0 .net "out", 0 0, L_0x5c7c33120440;  alias, 1 drivers
S_0x5c7c32e937a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e93580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120440 .functor NAND 1, L_0x5c7c33120390, L_0x5c7c33120390, C4<1>, C4<1>;
v0x5c7c32e93a10_0 .net "in_a", 0 0, L_0x5c7c33120390;  alias, 1 drivers
v0x5c7c32e93ad0_0 .net "in_b", 0 0, L_0x5c7c33120390;  alias, 1 drivers
v0x5c7c32e93c20_0 .net "out", 0 0, L_0x5c7c33120440;  alias, 1 drivers
S_0x5c7c32e94fa0 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32e7ce30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e9a990_0 .net "branch1_out", 0 0, L_0x5c7c331206d0;  1 drivers
v0x5c7c32e9aac0_0 .net "branch2_out", 0 0, L_0x5c7c33120960;  1 drivers
v0x5c7c32e9ac10_0 .net "in_a", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e9adf0_0 .net "in_b", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e9afa0_0 .net "out", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32e9b040_0 .net "temp1_out", 0 0, L_0x5c7c33120620;  1 drivers
v0x5c7c32e9b0e0_0 .net "temp2_out", 0 0, L_0x5c7c331208b0;  1 drivers
v0x5c7c32e9b180_0 .net "temp3_out", 0 0, L_0x5c7c33120b40;  1 drivers
S_0x5c7c32e95130 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32e94fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e961d0_0 .net "in_a", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e96270_0 .net "in_b", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e96330_0 .net "out", 0 0, L_0x5c7c33120620;  alias, 1 drivers
v0x5c7c32e96450_0 .net "temp_out", 0 0, L_0x5c7c32e93bb0;  1 drivers
S_0x5c7c32e95350 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e95130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e93bb0 .functor NAND 1, L_0x5c7c3311e9c0, L_0x5c7c3311e9c0, C4<1>, C4<1>;
v0x5c7c32e955c0_0 .net "in_a", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e95710_0 .net "in_b", 0 0, L_0x5c7c3311e9c0;  alias, 1 drivers
v0x5c7c32e957d0_0 .net "out", 0 0, L_0x5c7c32e93bb0;  alias, 1 drivers
S_0x5c7c32e95900 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e95130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e96020_0 .net "in_a", 0 0, L_0x5c7c32e93bb0;  alias, 1 drivers
v0x5c7c32e960c0_0 .net "out", 0 0, L_0x5c7c33120620;  alias, 1 drivers
S_0x5c7c32e95ad0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e95900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120620 .functor NAND 1, L_0x5c7c32e93bb0, L_0x5c7c32e93bb0, C4<1>, C4<1>;
v0x5c7c32e95d40_0 .net "in_a", 0 0, L_0x5c7c32e93bb0;  alias, 1 drivers
v0x5c7c32e95e30_0 .net "in_b", 0 0, L_0x5c7c32e93bb0;  alias, 1 drivers
v0x5c7c32e95f20_0 .net "out", 0 0, L_0x5c7c33120620;  alias, 1 drivers
S_0x5c7c32e965c0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32e94fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e975f0_0 .net "in_a", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e97690_0 .net "in_b", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e97750_0 .net "out", 0 0, L_0x5c7c331208b0;  alias, 1 drivers
v0x5c7c32e97870_0 .net "temp_out", 0 0, L_0x5c7c32e99410;  1 drivers
S_0x5c7c32e967a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e965c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e99410 .functor NAND 1, L_0x5c7c3311fb10, L_0x5c7c3311fb10, C4<1>, C4<1>;
v0x5c7c32e96a10_0 .net "in_a", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e96b60_0 .net "in_b", 0 0, L_0x5c7c3311fb10;  alias, 1 drivers
v0x5c7c32e96c20_0 .net "out", 0 0, L_0x5c7c32e99410;  alias, 1 drivers
S_0x5c7c32e96d20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e965c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e97440_0 .net "in_a", 0 0, L_0x5c7c32e99410;  alias, 1 drivers
v0x5c7c32e974e0_0 .net "out", 0 0, L_0x5c7c331208b0;  alias, 1 drivers
S_0x5c7c32e96ef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e96d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331208b0 .functor NAND 1, L_0x5c7c32e99410, L_0x5c7c32e99410, C4<1>, C4<1>;
v0x5c7c32e97160_0 .net "in_a", 0 0, L_0x5c7c32e99410;  alias, 1 drivers
v0x5c7c32e97250_0 .net "in_b", 0 0, L_0x5c7c32e99410;  alias, 1 drivers
v0x5c7c32e97340_0 .net "out", 0 0, L_0x5c7c331208b0;  alias, 1 drivers
S_0x5c7c32e979e0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32e94fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e98a20_0 .net "in_a", 0 0, L_0x5c7c331206d0;  alias, 1 drivers
v0x5c7c32e98af0_0 .net "in_b", 0 0, L_0x5c7c33120960;  alias, 1 drivers
v0x5c7c32e98bc0_0 .net "out", 0 0, L_0x5c7c33120b40;  alias, 1 drivers
v0x5c7c32e98ce0_0 .net "temp_out", 0 0, L_0x5c7c32e99d80;  1 drivers
S_0x5c7c32e97bc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e979e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e99d80 .functor NAND 1, L_0x5c7c331206d0, L_0x5c7c33120960, C4<1>, C4<1>;
v0x5c7c32e97e10_0 .net "in_a", 0 0, L_0x5c7c331206d0;  alias, 1 drivers
v0x5c7c32e97ef0_0 .net "in_b", 0 0, L_0x5c7c33120960;  alias, 1 drivers
v0x5c7c32e97fb0_0 .net "out", 0 0, L_0x5c7c32e99d80;  alias, 1 drivers
S_0x5c7c32e98100 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e979e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e98870_0 .net "in_a", 0 0, L_0x5c7c32e99d80;  alias, 1 drivers
v0x5c7c32e98910_0 .net "out", 0 0, L_0x5c7c33120b40;  alias, 1 drivers
S_0x5c7c32e98320 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e98100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120b40 .functor NAND 1, L_0x5c7c32e99d80, L_0x5c7c32e99d80, C4<1>, C4<1>;
v0x5c7c32e98590_0 .net "in_a", 0 0, L_0x5c7c32e99d80;  alias, 1 drivers
v0x5c7c32e98680_0 .net "in_b", 0 0, L_0x5c7c32e99d80;  alias, 1 drivers
v0x5c7c32e98770_0 .net "out", 0 0, L_0x5c7c33120b40;  alias, 1 drivers
S_0x5c7c32e98e30 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32e94fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e99560_0 .net "in_a", 0 0, L_0x5c7c33120620;  alias, 1 drivers
v0x5c7c32e99600_0 .net "out", 0 0, L_0x5c7c331206d0;  alias, 1 drivers
S_0x5c7c32e99000 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e98e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331206d0 .functor NAND 1, L_0x5c7c33120620, L_0x5c7c33120620, C4<1>, C4<1>;
v0x5c7c32e99270_0 .net "in_a", 0 0, L_0x5c7c33120620;  alias, 1 drivers
v0x5c7c32e99330_0 .net "in_b", 0 0, L_0x5c7c33120620;  alias, 1 drivers
v0x5c7c32e99480_0 .net "out", 0 0, L_0x5c7c331206d0;  alias, 1 drivers
S_0x5c7c32e99700 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32e94fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e99ed0_0 .net "in_a", 0 0, L_0x5c7c331208b0;  alias, 1 drivers
v0x5c7c32e99f70_0 .net "out", 0 0, L_0x5c7c33120960;  alias, 1 drivers
S_0x5c7c32e99970 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e99700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120960 .functor NAND 1, L_0x5c7c331208b0, L_0x5c7c331208b0, C4<1>, C4<1>;
v0x5c7c32e99be0_0 .net "in_a", 0 0, L_0x5c7c331208b0;  alias, 1 drivers
v0x5c7c32e99ca0_0 .net "in_b", 0 0, L_0x5c7c331208b0;  alias, 1 drivers
v0x5c7c32e99df0_0 .net "out", 0 0, L_0x5c7c33120960;  alias, 1 drivers
S_0x5c7c32e9a070 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32e94fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e9a810_0 .net "in_a", 0 0, L_0x5c7c33120b40;  alias, 1 drivers
v0x5c7c32e9a8b0_0 .net "out", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
S_0x5c7c32e9a290 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e9a070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120bf0 .functor NAND 1, L_0x5c7c33120b40, L_0x5c7c33120b40, C4<1>, C4<1>;
v0x5c7c32e9a500_0 .net "in_a", 0 0, L_0x5c7c33120b40;  alias, 1 drivers
v0x5c7c32e9a5c0_0 .net "in_b", 0 0, L_0x5c7c33120b40;  alias, 1 drivers
v0x5c7c32e9a710_0 .net "out", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
S_0x5c7c32e9b7e0 .scope module, "fa_gate8" "FullAdder" 2 13, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32ed9c10_0 .net "a", 0 0, L_0x5c7c33123300;  1 drivers
v0x5c7c32ed9cb0_0 .net "b", 0 0, L_0x5c7c331234b0;  1 drivers
v0x5c7c32ed9d70_0 .net "c", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ed9e10_0 .net "carry", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ed9eb0_0 .net "sum", 0 0, L_0x5c7c331229b0;  1 drivers
v0x5c7c32ed9f50_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33120f50;  1 drivers
v0x5c7c32ed9ff0_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33122080;  1 drivers
v0x5c7c32eda090_0 .net "tmp_sum_out", 0 0, L_0x5c7c33121a80;  1 drivers
S_0x5c7c32e9ba40 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32e9b7e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32ea75c0_0 .net "a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32ea7770_0 .net "b", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32ea7940_0 .net "carry", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32ea79e0_0 .net "sum", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
S_0x5c7c32e9bcb0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32e9ba40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e9cda0_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32e9ce70_0 .net "in_b", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32e9cf40_0 .net "out", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32e9d060_0 .net "temp_out", 0 0, L_0x5c7c32e5d340;  1 drivers
S_0x5c7c32e9bf20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e9bcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32e5d340 .functor NAND 1, L_0x5c7c33123300, L_0x5c7c331234b0, C4<1>, C4<1>;
v0x5c7c32e9c190_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32e9c270_0 .net "in_b", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32e9c330_0 .net "out", 0 0, L_0x5c7c32e5d340;  alias, 1 drivers
S_0x5c7c32e9c480 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e9bcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e9cbf0_0 .net "in_a", 0 0, L_0x5c7c32e5d340;  alias, 1 drivers
v0x5c7c32e9cc90_0 .net "out", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
S_0x5c7c32e9c6a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e9c480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120f50 .functor NAND 1, L_0x5c7c32e5d340, L_0x5c7c32e5d340, C4<1>, C4<1>;
v0x5c7c32e9c910_0 .net "in_a", 0 0, L_0x5c7c32e5d340;  alias, 1 drivers
v0x5c7c32e9ca00_0 .net "in_b", 0 0, L_0x5c7c32e5d340;  alias, 1 drivers
v0x5c7c32e9caf0_0 .net "out", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
S_0x5c7c32e9d120 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32e9ba40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ea6ee0_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32ea6f80_0 .net "in_b", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32ea7040_0 .net "out", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ea70e0_0 .net "temp_a_and_out", 0 0, L_0x5c7c33121140;  1 drivers
v0x5c7c32ea7290_0 .net "temp_a_out", 0 0, L_0x5c7c33120fe0;  1 drivers
v0x5c7c32ea7330_0 .net "temp_b_and_out", 0 0, L_0x5c7c33121350;  1 drivers
v0x5c7c32ea74e0_0 .net "temp_b_out", 0 0, L_0x5c7c331211f0;  1 drivers
S_0x5c7c32e9d300 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32e9d120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e9e3c0_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32e9e460_0 .net "in_b", 0 0, L_0x5c7c33120fe0;  alias, 1 drivers
v0x5c7c32e9e550_0 .net "out", 0 0, L_0x5c7c33121140;  alias, 1 drivers
v0x5c7c32e9e670_0 .net "temp_out", 0 0, L_0x5c7c33121090;  1 drivers
S_0x5c7c32e9d570 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e9d300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121090 .functor NAND 1, L_0x5c7c33123300, L_0x5c7c33120fe0, C4<1>, C4<1>;
v0x5c7c32e9d7e0_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32e9d8f0_0 .net "in_b", 0 0, L_0x5c7c33120fe0;  alias, 1 drivers
v0x5c7c32e9d9b0_0 .net "out", 0 0, L_0x5c7c33121090;  alias, 1 drivers
S_0x5c7c32e9dad0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e9d300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e9e210_0 .net "in_a", 0 0, L_0x5c7c33121090;  alias, 1 drivers
v0x5c7c32e9e2b0_0 .net "out", 0 0, L_0x5c7c33121140;  alias, 1 drivers
S_0x5c7c32e9dcf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e9dad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121140 .functor NAND 1, L_0x5c7c33121090, L_0x5c7c33121090, C4<1>, C4<1>;
v0x5c7c32e9df60_0 .net "in_a", 0 0, L_0x5c7c33121090;  alias, 1 drivers
v0x5c7c32e9e020_0 .net "in_b", 0 0, L_0x5c7c33121090;  alias, 1 drivers
v0x5c7c32e9e110_0 .net "out", 0 0, L_0x5c7c33121140;  alias, 1 drivers
S_0x5c7c32e9e730 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32e9d120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32e9f760_0 .net "in_a", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32e9f800_0 .net "in_b", 0 0, L_0x5c7c331211f0;  alias, 1 drivers
v0x5c7c32e9f8f0_0 .net "out", 0 0, L_0x5c7c33121350;  alias, 1 drivers
v0x5c7c32e9fa10_0 .net "temp_out", 0 0, L_0x5c7c331212a0;  1 drivers
S_0x5c7c32e9e910 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32e9e730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331212a0 .functor NAND 1, L_0x5c7c331234b0, L_0x5c7c331211f0, C4<1>, C4<1>;
v0x5c7c32e9eb80_0 .net "in_a", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32e9ec90_0 .net "in_b", 0 0, L_0x5c7c331211f0;  alias, 1 drivers
v0x5c7c32e9ed50_0 .net "out", 0 0, L_0x5c7c331212a0;  alias, 1 drivers
S_0x5c7c32e9ee70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32e9e730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32e9f5b0_0 .net "in_a", 0 0, L_0x5c7c331212a0;  alias, 1 drivers
v0x5c7c32e9f650_0 .net "out", 0 0, L_0x5c7c33121350;  alias, 1 drivers
S_0x5c7c32e9f090 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e9ee70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121350 .functor NAND 1, L_0x5c7c331212a0, L_0x5c7c331212a0, C4<1>, C4<1>;
v0x5c7c32e9f300_0 .net "in_a", 0 0, L_0x5c7c331212a0;  alias, 1 drivers
v0x5c7c32e9f3c0_0 .net "in_b", 0 0, L_0x5c7c331212a0;  alias, 1 drivers
v0x5c7c32e9f4b0_0 .net "out", 0 0, L_0x5c7c33121350;  alias, 1 drivers
S_0x5c7c32e9fb60 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32e9d120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea02a0_0 .net "in_a", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32ea0340_0 .net "out", 0 0, L_0x5c7c33120fe0;  alias, 1 drivers
S_0x5c7c32e9fd30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32e9fb60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33120fe0 .functor NAND 1, L_0x5c7c331234b0, L_0x5c7c331234b0, C4<1>, C4<1>;
v0x5c7c32e9ff80_0 .net "in_a", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32ea00d0_0 .net "in_b", 0 0, L_0x5c7c331234b0;  alias, 1 drivers
v0x5c7c32ea0190_0 .net "out", 0 0, L_0x5c7c33120fe0;  alias, 1 drivers
S_0x5c7c32ea0440 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32e9d120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea0bc0_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32ea0c60_0 .net "out", 0 0, L_0x5c7c331211f0;  alias, 1 drivers
S_0x5c7c32ea0660 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea0440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331211f0 .functor NAND 1, L_0x5c7c33123300, L_0x5c7c33123300, C4<1>, C4<1>;
v0x5c7c32ea08d0_0 .net "in_a", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32ea0a20_0 .net "in_b", 0 0, L_0x5c7c33123300;  alias, 1 drivers
v0x5c7c32ea0ae0_0 .net "out", 0 0, L_0x5c7c331211f0;  alias, 1 drivers
S_0x5c7c32ea0d60 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32e9d120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ea6830_0 .net "branch1_out", 0 0, L_0x5c7c33121560;  1 drivers
v0x5c7c32ea6960_0 .net "branch2_out", 0 0, L_0x5c7c331217f0;  1 drivers
v0x5c7c32ea6ab0_0 .net "in_a", 0 0, L_0x5c7c33121140;  alias, 1 drivers
v0x5c7c32ea6b80_0 .net "in_b", 0 0, L_0x5c7c33121350;  alias, 1 drivers
v0x5c7c32ea6c20_0 .net "out", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ea6cc0_0 .net "temp1_out", 0 0, L_0x5c7c331214b0;  1 drivers
v0x5c7c32ea6d60_0 .net "temp2_out", 0 0, L_0x5c7c33121740;  1 drivers
v0x5c7c32ea6e00_0 .net "temp3_out", 0 0, L_0x5c7c331219d0;  1 drivers
S_0x5c7c32ea0fe0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32ea0d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ea2070_0 .net "in_a", 0 0, L_0x5c7c33121140;  alias, 1 drivers
v0x5c7c32ea2110_0 .net "in_b", 0 0, L_0x5c7c33121140;  alias, 1 drivers
v0x5c7c32ea21d0_0 .net "out", 0 0, L_0x5c7c331214b0;  alias, 1 drivers
v0x5c7c32ea22f0_0 .net "temp_out", 0 0, L_0x5c7c33121400;  1 drivers
S_0x5c7c32ea1250 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ea0fe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121400 .functor NAND 1, L_0x5c7c33121140, L_0x5c7c33121140, C4<1>, C4<1>;
v0x5c7c32ea14c0_0 .net "in_a", 0 0, L_0x5c7c33121140;  alias, 1 drivers
v0x5c7c32ea1580_0 .net "in_b", 0 0, L_0x5c7c33121140;  alias, 1 drivers
v0x5c7c32ea16d0_0 .net "out", 0 0, L_0x5c7c33121400;  alias, 1 drivers
S_0x5c7c32ea17d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ea0fe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea1ec0_0 .net "in_a", 0 0, L_0x5c7c33121400;  alias, 1 drivers
v0x5c7c32ea1f60_0 .net "out", 0 0, L_0x5c7c331214b0;  alias, 1 drivers
S_0x5c7c32ea19a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea17d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331214b0 .functor NAND 1, L_0x5c7c33121400, L_0x5c7c33121400, C4<1>, C4<1>;
v0x5c7c32ea1c10_0 .net "in_a", 0 0, L_0x5c7c33121400;  alias, 1 drivers
v0x5c7c32ea1cd0_0 .net "in_b", 0 0, L_0x5c7c33121400;  alias, 1 drivers
v0x5c7c32ea1dc0_0 .net "out", 0 0, L_0x5c7c331214b0;  alias, 1 drivers
S_0x5c7c32ea2460 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32ea0d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ea3490_0 .net "in_a", 0 0, L_0x5c7c33121350;  alias, 1 drivers
v0x5c7c32ea3530_0 .net "in_b", 0 0, L_0x5c7c33121350;  alias, 1 drivers
v0x5c7c32ea35f0_0 .net "out", 0 0, L_0x5c7c33121740;  alias, 1 drivers
v0x5c7c32ea3710_0 .net "temp_out", 0 0, L_0x5c7c32ea52b0;  1 drivers
S_0x5c7c32ea2640 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ea2460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ea52b0 .functor NAND 1, L_0x5c7c33121350, L_0x5c7c33121350, C4<1>, C4<1>;
v0x5c7c32ea28b0_0 .net "in_a", 0 0, L_0x5c7c33121350;  alias, 1 drivers
v0x5c7c32ea2970_0 .net "in_b", 0 0, L_0x5c7c33121350;  alias, 1 drivers
v0x5c7c32ea2ac0_0 .net "out", 0 0, L_0x5c7c32ea52b0;  alias, 1 drivers
S_0x5c7c32ea2bc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ea2460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea32e0_0 .net "in_a", 0 0, L_0x5c7c32ea52b0;  alias, 1 drivers
v0x5c7c32ea3380_0 .net "out", 0 0, L_0x5c7c33121740;  alias, 1 drivers
S_0x5c7c32ea2d90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea2bc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121740 .functor NAND 1, L_0x5c7c32ea52b0, L_0x5c7c32ea52b0, C4<1>, C4<1>;
v0x5c7c32ea3000_0 .net "in_a", 0 0, L_0x5c7c32ea52b0;  alias, 1 drivers
v0x5c7c32ea30f0_0 .net "in_b", 0 0, L_0x5c7c32ea52b0;  alias, 1 drivers
v0x5c7c32ea31e0_0 .net "out", 0 0, L_0x5c7c33121740;  alias, 1 drivers
S_0x5c7c32ea3880 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32ea0d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ea48c0_0 .net "in_a", 0 0, L_0x5c7c33121560;  alias, 1 drivers
v0x5c7c32ea4990_0 .net "in_b", 0 0, L_0x5c7c331217f0;  alias, 1 drivers
v0x5c7c32ea4a60_0 .net "out", 0 0, L_0x5c7c331219d0;  alias, 1 drivers
v0x5c7c32ea4b80_0 .net "temp_out", 0 0, L_0x5c7c32ea5c20;  1 drivers
S_0x5c7c32ea3a60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ea3880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ea5c20 .functor NAND 1, L_0x5c7c33121560, L_0x5c7c331217f0, C4<1>, C4<1>;
v0x5c7c32ea3cb0_0 .net "in_a", 0 0, L_0x5c7c33121560;  alias, 1 drivers
v0x5c7c32ea3d90_0 .net "in_b", 0 0, L_0x5c7c331217f0;  alias, 1 drivers
v0x5c7c32ea3e50_0 .net "out", 0 0, L_0x5c7c32ea5c20;  alias, 1 drivers
S_0x5c7c32ea3fa0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ea3880;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea4710_0 .net "in_a", 0 0, L_0x5c7c32ea5c20;  alias, 1 drivers
v0x5c7c32ea47b0_0 .net "out", 0 0, L_0x5c7c331219d0;  alias, 1 drivers
S_0x5c7c32ea41c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea3fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331219d0 .functor NAND 1, L_0x5c7c32ea5c20, L_0x5c7c32ea5c20, C4<1>, C4<1>;
v0x5c7c32ea4430_0 .net "in_a", 0 0, L_0x5c7c32ea5c20;  alias, 1 drivers
v0x5c7c32ea4520_0 .net "in_b", 0 0, L_0x5c7c32ea5c20;  alias, 1 drivers
v0x5c7c32ea4610_0 .net "out", 0 0, L_0x5c7c331219d0;  alias, 1 drivers
S_0x5c7c32ea4cd0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32ea0d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea5400_0 .net "in_a", 0 0, L_0x5c7c331214b0;  alias, 1 drivers
v0x5c7c32ea54a0_0 .net "out", 0 0, L_0x5c7c33121560;  alias, 1 drivers
S_0x5c7c32ea4ea0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea4cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121560 .functor NAND 1, L_0x5c7c331214b0, L_0x5c7c331214b0, C4<1>, C4<1>;
v0x5c7c32ea5110_0 .net "in_a", 0 0, L_0x5c7c331214b0;  alias, 1 drivers
v0x5c7c32ea51d0_0 .net "in_b", 0 0, L_0x5c7c331214b0;  alias, 1 drivers
v0x5c7c32ea5320_0 .net "out", 0 0, L_0x5c7c33121560;  alias, 1 drivers
S_0x5c7c32ea55a0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32ea0d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea5d70_0 .net "in_a", 0 0, L_0x5c7c33121740;  alias, 1 drivers
v0x5c7c32ea5e10_0 .net "out", 0 0, L_0x5c7c331217f0;  alias, 1 drivers
S_0x5c7c32ea5810 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea55a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331217f0 .functor NAND 1, L_0x5c7c33121740, L_0x5c7c33121740, C4<1>, C4<1>;
v0x5c7c32ea5a80_0 .net "in_a", 0 0, L_0x5c7c33121740;  alias, 1 drivers
v0x5c7c32ea5b40_0 .net "in_b", 0 0, L_0x5c7c33121740;  alias, 1 drivers
v0x5c7c32ea5c90_0 .net "out", 0 0, L_0x5c7c331217f0;  alias, 1 drivers
S_0x5c7c32ea5f10 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32ea0d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea66b0_0 .net "in_a", 0 0, L_0x5c7c331219d0;  alias, 1 drivers
v0x5c7c32ea6750_0 .net "out", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
S_0x5c7c32ea6130 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea5f10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33121a80 .functor NAND 1, L_0x5c7c331219d0, L_0x5c7c331219d0, C4<1>, C4<1>;
v0x5c7c32ea63a0_0 .net "in_a", 0 0, L_0x5c7c331219d0;  alias, 1 drivers
v0x5c7c32ea6460_0 .net "in_b", 0 0, L_0x5c7c331219d0;  alias, 1 drivers
v0x5c7c32ea65b0_0 .net "out", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
S_0x5c7c32ea7ac0 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32e9b7e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32ed35e0_0 .net "a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ed3680_0 .net "b", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ed3740_0 .net "carry", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ed37e0_0 .net "sum", 0 0, L_0x5c7c331229b0;  alias, 1 drivers
S_0x5c7c32ea7ce0 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32ea7ac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ea8c80_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ea8d20_0 .net "in_b", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ea8de0_0 .net "out", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ea8f00_0 .net "temp_out", 0 0, L_0x5c7c32ea6540;  1 drivers
S_0x5c7c32ea7e90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ea7ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ea6540 .functor NAND 1, L_0x5c7c33121a80, L_0x5c7c33120bf0, C4<1>, C4<1>;
v0x5c7c32ea8100_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ea81c0_0 .net "in_b", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ea8280_0 .net "out", 0 0, L_0x5c7c32ea6540;  alias, 1 drivers
S_0x5c7c32ea83b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ea7ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ea8ad0_0 .net "in_a", 0 0, L_0x5c7c32ea6540;  alias, 1 drivers
v0x5c7c32ea8b70_0 .net "out", 0 0, L_0x5c7c33122080;  alias, 1 drivers
S_0x5c7c32ea8580 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea83b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122080 .functor NAND 1, L_0x5c7c32ea6540, L_0x5c7c32ea6540, C4<1>, C4<1>;
v0x5c7c32ea87f0_0 .net "in_a", 0 0, L_0x5c7c32ea6540;  alias, 1 drivers
v0x5c7c32ea88e0_0 .net "in_b", 0 0, L_0x5c7c32ea6540;  alias, 1 drivers
v0x5c7c32ea89d0_0 .net "out", 0 0, L_0x5c7c33122080;  alias, 1 drivers
S_0x5c7c32ea9070 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32ea7ac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed2f00_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ed2fa0_0 .net "in_b", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ed3060_0 .net "out", 0 0, L_0x5c7c331229b0;  alias, 1 drivers
v0x5c7c32ed3100_0 .net "temp_a_and_out", 0 0, L_0x5c7c33122290;  1 drivers
v0x5c7c32ed32b0_0 .net "temp_a_out", 0 0, L_0x5c7c33122130;  1 drivers
v0x5c7c32ed3350_0 .net "temp_b_and_out", 0 0, L_0x5c7c331224a0;  1 drivers
v0x5c7c32ed3500_0 .net "temp_b_out", 0 0, L_0x5c7c33122340;  1 drivers
S_0x5c7c32ea9250 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32ea9070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32eaa2f0_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32eaa4a0_0 .net "in_b", 0 0, L_0x5c7c33122130;  alias, 1 drivers
v0x5c7c32eaa590_0 .net "out", 0 0, L_0x5c7c33122290;  alias, 1 drivers
v0x5c7c32eaa6b0_0 .net "temp_out", 0 0, L_0x5c7c331221e0;  1 drivers
S_0x5c7c32ea94c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ea9250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331221e0 .functor NAND 1, L_0x5c7c33121a80, L_0x5c7c33122130, C4<1>, C4<1>;
v0x5c7c32ea9730_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ea97f0_0 .net "in_b", 0 0, L_0x5c7c33122130;  alias, 1 drivers
v0x5c7c32ea98b0_0 .net "out", 0 0, L_0x5c7c331221e0;  alias, 1 drivers
S_0x5c7c32ea99d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ea9250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eaa140_0 .net "in_a", 0 0, L_0x5c7c331221e0;  alias, 1 drivers
v0x5c7c32eaa1e0_0 .net "out", 0 0, L_0x5c7c33122290;  alias, 1 drivers
S_0x5c7c32ea9bf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ea99d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122290 .functor NAND 1, L_0x5c7c331221e0, L_0x5c7c331221e0, C4<1>, C4<1>;
v0x5c7c32ea9e60_0 .net "in_a", 0 0, L_0x5c7c331221e0;  alias, 1 drivers
v0x5c7c32ea9f50_0 .net "in_b", 0 0, L_0x5c7c331221e0;  alias, 1 drivers
v0x5c7c32eaa040_0 .net "out", 0 0, L_0x5c7c33122290;  alias, 1 drivers
S_0x5c7c32eaa770 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32ea9070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ecb780_0 .net "in_a", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ecb820_0 .net "in_b", 0 0, L_0x5c7c33122340;  alias, 1 drivers
v0x5c7c32ecb910_0 .net "out", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
v0x5c7c32ecba30_0 .net "temp_out", 0 0, L_0x5c7c331223f0;  1 drivers
S_0x5c7c32eaa950 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32eaa770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331223f0 .functor NAND 1, L_0x5c7c33120bf0, L_0x5c7c33122340, C4<1>, C4<1>;
v0x5c7c32eaabc0_0 .net "in_a", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32eaac80_0 .net "in_b", 0 0, L_0x5c7c33122340;  alias, 1 drivers
v0x5c7c32eaad40_0 .net "out", 0 0, L_0x5c7c331223f0;  alias, 1 drivers
S_0x5c7c32eaae60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32eaa770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ecb5d0_0 .net "in_a", 0 0, L_0x5c7c331223f0;  alias, 1 drivers
v0x5c7c32ecb670_0 .net "out", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
S_0x5c7c32eab080 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eaae60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331224a0 .functor NAND 1, L_0x5c7c331223f0, L_0x5c7c331223f0, C4<1>, C4<1>;
v0x5c7c32eab2f0_0 .net "in_a", 0 0, L_0x5c7c331223f0;  alias, 1 drivers
v0x5c7c32eab3e0_0 .net "in_b", 0 0, L_0x5c7c331223f0;  alias, 1 drivers
v0x5c7c32eab4d0_0 .net "out", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
S_0x5c7c32ecbb80 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32ea9070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ecc390_0 .net "in_a", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ecc430_0 .net "out", 0 0, L_0x5c7c33122130;  alias, 1 drivers
S_0x5c7c32ecbd50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ecbb80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122130 .functor NAND 1, L_0x5c7c33120bf0, L_0x5c7c33120bf0, C4<1>, C4<1>;
v0x5c7c32ecbfa0_0 .net "in_a", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ecc170_0 .net "in_b", 0 0, L_0x5c7c33120bf0;  alias, 1 drivers
v0x5c7c32ecc230_0 .net "out", 0 0, L_0x5c7c33122130;  alias, 1 drivers
S_0x5c7c32ecc530 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32ea9070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eccc70_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32eccd10_0 .net "out", 0 0, L_0x5c7c33122340;  alias, 1 drivers
S_0x5c7c32ecc750 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ecc530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122340 .functor NAND 1, L_0x5c7c33121a80, L_0x5c7c33121a80, C4<1>, C4<1>;
v0x5c7c32ecc9c0_0 .net "in_a", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32ecca80_0 .net "in_b", 0 0, L_0x5c7c33121a80;  alias, 1 drivers
v0x5c7c32eccb40_0 .net "out", 0 0, L_0x5c7c33122340;  alias, 1 drivers
S_0x5c7c32ecce10 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32ea9070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed2850_0 .net "branch1_out", 0 0, L_0x5c7c331226b0;  1 drivers
v0x5c7c32ed2980_0 .net "branch2_out", 0 0, L_0x5c7c33122830;  1 drivers
v0x5c7c32ed2ad0_0 .net "in_a", 0 0, L_0x5c7c33122290;  alias, 1 drivers
v0x5c7c32ed2ba0_0 .net "in_b", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
v0x5c7c32ed2c40_0 .net "out", 0 0, L_0x5c7c331229b0;  alias, 1 drivers
v0x5c7c32ed2ce0_0 .net "temp1_out", 0 0, L_0x5c7c33122600;  1 drivers
v0x5c7c32ed2d80_0 .net "temp2_out", 0 0, L_0x5c7c33122780;  1 drivers
v0x5c7c32ed2e20_0 .net "temp3_out", 0 0, L_0x5c7c33122900;  1 drivers
S_0x5c7c32ecd090 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32ecce10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ece090_0 .net "in_a", 0 0, L_0x5c7c33122290;  alias, 1 drivers
v0x5c7c32ece130_0 .net "in_b", 0 0, L_0x5c7c33122290;  alias, 1 drivers
v0x5c7c32ece1f0_0 .net "out", 0 0, L_0x5c7c33122600;  alias, 1 drivers
v0x5c7c32ece310_0 .net "temp_out", 0 0, L_0x5c7c33122550;  1 drivers
S_0x5c7c32ecd300 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ecd090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122550 .functor NAND 1, L_0x5c7c33122290, L_0x5c7c33122290, C4<1>, C4<1>;
v0x5c7c32ecd570_0 .net "in_a", 0 0, L_0x5c7c33122290;  alias, 1 drivers
v0x5c7c32ecd630_0 .net "in_b", 0 0, L_0x5c7c33122290;  alias, 1 drivers
v0x5c7c32ecd6f0_0 .net "out", 0 0, L_0x5c7c33122550;  alias, 1 drivers
S_0x5c7c32ecd7f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ecd090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ecdee0_0 .net "in_a", 0 0, L_0x5c7c33122550;  alias, 1 drivers
v0x5c7c32ecdf80_0 .net "out", 0 0, L_0x5c7c33122600;  alias, 1 drivers
S_0x5c7c32ecd9c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ecd7f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122600 .functor NAND 1, L_0x5c7c33122550, L_0x5c7c33122550, C4<1>, C4<1>;
v0x5c7c32ecdc30_0 .net "in_a", 0 0, L_0x5c7c33122550;  alias, 1 drivers
v0x5c7c32ecdcf0_0 .net "in_b", 0 0, L_0x5c7c33122550;  alias, 1 drivers
v0x5c7c32ecdde0_0 .net "out", 0 0, L_0x5c7c33122600;  alias, 1 drivers
S_0x5c7c32ece480 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32ecce10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ecf4b0_0 .net "in_a", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
v0x5c7c32ecf550_0 .net "in_b", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
v0x5c7c32ecf610_0 .net "out", 0 0, L_0x5c7c33122780;  alias, 1 drivers
v0x5c7c32ecf730_0 .net "temp_out", 0 0, L_0x5c7c32ed12d0;  1 drivers
S_0x5c7c32ece660 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ece480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ed12d0 .functor NAND 1, L_0x5c7c331224a0, L_0x5c7c331224a0, C4<1>, C4<1>;
v0x5c7c32ece8d0_0 .net "in_a", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
v0x5c7c32ece990_0 .net "in_b", 0 0, L_0x5c7c331224a0;  alias, 1 drivers
v0x5c7c32eceae0_0 .net "out", 0 0, L_0x5c7c32ed12d0;  alias, 1 drivers
S_0x5c7c32ecebe0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ece480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ecf300_0 .net "in_a", 0 0, L_0x5c7c32ed12d0;  alias, 1 drivers
v0x5c7c32ecf3a0_0 .net "out", 0 0, L_0x5c7c33122780;  alias, 1 drivers
S_0x5c7c32ecedb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ecebe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122780 .functor NAND 1, L_0x5c7c32ed12d0, L_0x5c7c32ed12d0, C4<1>, C4<1>;
v0x5c7c32ecf020_0 .net "in_a", 0 0, L_0x5c7c32ed12d0;  alias, 1 drivers
v0x5c7c32ecf110_0 .net "in_b", 0 0, L_0x5c7c32ed12d0;  alias, 1 drivers
v0x5c7c32ecf200_0 .net "out", 0 0, L_0x5c7c33122780;  alias, 1 drivers
S_0x5c7c32ecf8a0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32ecce10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed08e0_0 .net "in_a", 0 0, L_0x5c7c331226b0;  alias, 1 drivers
v0x5c7c32ed09b0_0 .net "in_b", 0 0, L_0x5c7c33122830;  alias, 1 drivers
v0x5c7c32ed0a80_0 .net "out", 0 0, L_0x5c7c33122900;  alias, 1 drivers
v0x5c7c32ed0ba0_0 .net "temp_out", 0 0, L_0x5c7c32ed1c40;  1 drivers
S_0x5c7c32ecfa80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ecf8a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ed1c40 .functor NAND 1, L_0x5c7c331226b0, L_0x5c7c33122830, C4<1>, C4<1>;
v0x5c7c32ecfcd0_0 .net "in_a", 0 0, L_0x5c7c331226b0;  alias, 1 drivers
v0x5c7c32ecfdb0_0 .net "in_b", 0 0, L_0x5c7c33122830;  alias, 1 drivers
v0x5c7c32ecfe70_0 .net "out", 0 0, L_0x5c7c32ed1c40;  alias, 1 drivers
S_0x5c7c32ecffc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ecf8a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed0730_0 .net "in_a", 0 0, L_0x5c7c32ed1c40;  alias, 1 drivers
v0x5c7c32ed07d0_0 .net "out", 0 0, L_0x5c7c33122900;  alias, 1 drivers
S_0x5c7c32ed01e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ecffc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122900 .functor NAND 1, L_0x5c7c32ed1c40, L_0x5c7c32ed1c40, C4<1>, C4<1>;
v0x5c7c32ed0450_0 .net "in_a", 0 0, L_0x5c7c32ed1c40;  alias, 1 drivers
v0x5c7c32ed0540_0 .net "in_b", 0 0, L_0x5c7c32ed1c40;  alias, 1 drivers
v0x5c7c32ed0630_0 .net "out", 0 0, L_0x5c7c33122900;  alias, 1 drivers
S_0x5c7c32ed0cf0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32ecce10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed1420_0 .net "in_a", 0 0, L_0x5c7c33122600;  alias, 1 drivers
v0x5c7c32ed14c0_0 .net "out", 0 0, L_0x5c7c331226b0;  alias, 1 drivers
S_0x5c7c32ed0ec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed0cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331226b0 .functor NAND 1, L_0x5c7c33122600, L_0x5c7c33122600, C4<1>, C4<1>;
v0x5c7c32ed1130_0 .net "in_a", 0 0, L_0x5c7c33122600;  alias, 1 drivers
v0x5c7c32ed11f0_0 .net "in_b", 0 0, L_0x5c7c33122600;  alias, 1 drivers
v0x5c7c32ed1340_0 .net "out", 0 0, L_0x5c7c331226b0;  alias, 1 drivers
S_0x5c7c32ed15c0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32ecce10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed1d90_0 .net "in_a", 0 0, L_0x5c7c33122780;  alias, 1 drivers
v0x5c7c32ed1e30_0 .net "out", 0 0, L_0x5c7c33122830;  alias, 1 drivers
S_0x5c7c32ed1830 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed15c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122830 .functor NAND 1, L_0x5c7c33122780, L_0x5c7c33122780, C4<1>, C4<1>;
v0x5c7c32ed1aa0_0 .net "in_a", 0 0, L_0x5c7c33122780;  alias, 1 drivers
v0x5c7c32ed1b60_0 .net "in_b", 0 0, L_0x5c7c33122780;  alias, 1 drivers
v0x5c7c32ed1cb0_0 .net "out", 0 0, L_0x5c7c33122830;  alias, 1 drivers
S_0x5c7c32ed1f30 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32ecce10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed26d0_0 .net "in_a", 0 0, L_0x5c7c33122900;  alias, 1 drivers
v0x5c7c32ed2770_0 .net "out", 0 0, L_0x5c7c331229b0;  alias, 1 drivers
S_0x5c7c32ed2150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed1f30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331229b0 .functor NAND 1, L_0x5c7c33122900, L_0x5c7c33122900, C4<1>, C4<1>;
v0x5c7c32ed23c0_0 .net "in_a", 0 0, L_0x5c7c33122900;  alias, 1 drivers
v0x5c7c32ed2480_0 .net "in_b", 0 0, L_0x5c7c33122900;  alias, 1 drivers
v0x5c7c32ed25d0_0 .net "out", 0 0, L_0x5c7c331229b0;  alias, 1 drivers
S_0x5c7c32ed3950 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32e9b7e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed9340_0 .net "branch1_out", 0 0, L_0x5c7c33122c40;  1 drivers
v0x5c7c32ed9470_0 .net "branch2_out", 0 0, L_0x5c7c33122ed0;  1 drivers
v0x5c7c32ed95c0_0 .net "in_a", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32ed97a0_0 .net "in_b", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ed9950_0 .net "out", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ed99f0_0 .net "temp1_out", 0 0, L_0x5c7c33122b90;  1 drivers
v0x5c7c32ed9a90_0 .net "temp2_out", 0 0, L_0x5c7c33122e20;  1 drivers
v0x5c7c32ed9b30_0 .net "temp3_out", 0 0, L_0x5c7c331230b0;  1 drivers
S_0x5c7c32ed3ae0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32ed3950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed4b80_0 .net "in_a", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32ed4c20_0 .net "in_b", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32ed4ce0_0 .net "out", 0 0, L_0x5c7c33122b90;  alias, 1 drivers
v0x5c7c32ed4e00_0 .net "temp_out", 0 0, L_0x5c7c32ed2560;  1 drivers
S_0x5c7c32ed3d00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ed3ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ed2560 .functor NAND 1, L_0x5c7c33120f50, L_0x5c7c33120f50, C4<1>, C4<1>;
v0x5c7c32ed3f70_0 .net "in_a", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32ed40c0_0 .net "in_b", 0 0, L_0x5c7c33120f50;  alias, 1 drivers
v0x5c7c32ed4180_0 .net "out", 0 0, L_0x5c7c32ed2560;  alias, 1 drivers
S_0x5c7c32ed42b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ed3ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed49d0_0 .net "in_a", 0 0, L_0x5c7c32ed2560;  alias, 1 drivers
v0x5c7c32ed4a70_0 .net "out", 0 0, L_0x5c7c33122b90;  alias, 1 drivers
S_0x5c7c32ed4480 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed42b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122b90 .functor NAND 1, L_0x5c7c32ed2560, L_0x5c7c32ed2560, C4<1>, C4<1>;
v0x5c7c32ed46f0_0 .net "in_a", 0 0, L_0x5c7c32ed2560;  alias, 1 drivers
v0x5c7c32ed47e0_0 .net "in_b", 0 0, L_0x5c7c32ed2560;  alias, 1 drivers
v0x5c7c32ed48d0_0 .net "out", 0 0, L_0x5c7c33122b90;  alias, 1 drivers
S_0x5c7c32ed4f70 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32ed3950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed5fa0_0 .net "in_a", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ed6040_0 .net "in_b", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ed6100_0 .net "out", 0 0, L_0x5c7c33122e20;  alias, 1 drivers
v0x5c7c32ed6220_0 .net "temp_out", 0 0, L_0x5c7c32ed7dc0;  1 drivers
S_0x5c7c32ed5150 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ed4f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ed7dc0 .functor NAND 1, L_0x5c7c33122080, L_0x5c7c33122080, C4<1>, C4<1>;
v0x5c7c32ed53c0_0 .net "in_a", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ed5510_0 .net "in_b", 0 0, L_0x5c7c33122080;  alias, 1 drivers
v0x5c7c32ed55d0_0 .net "out", 0 0, L_0x5c7c32ed7dc0;  alias, 1 drivers
S_0x5c7c32ed56d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ed4f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed5df0_0 .net "in_a", 0 0, L_0x5c7c32ed7dc0;  alias, 1 drivers
v0x5c7c32ed5e90_0 .net "out", 0 0, L_0x5c7c33122e20;  alias, 1 drivers
S_0x5c7c32ed58a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed56d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122e20 .functor NAND 1, L_0x5c7c32ed7dc0, L_0x5c7c32ed7dc0, C4<1>, C4<1>;
v0x5c7c32ed5b10_0 .net "in_a", 0 0, L_0x5c7c32ed7dc0;  alias, 1 drivers
v0x5c7c32ed5c00_0 .net "in_b", 0 0, L_0x5c7c32ed7dc0;  alias, 1 drivers
v0x5c7c32ed5cf0_0 .net "out", 0 0, L_0x5c7c33122e20;  alias, 1 drivers
S_0x5c7c32ed6390 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32ed3950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ed73d0_0 .net "in_a", 0 0, L_0x5c7c33122c40;  alias, 1 drivers
v0x5c7c32ed74a0_0 .net "in_b", 0 0, L_0x5c7c33122ed0;  alias, 1 drivers
v0x5c7c32ed7570_0 .net "out", 0 0, L_0x5c7c331230b0;  alias, 1 drivers
v0x5c7c32ed7690_0 .net "temp_out", 0 0, L_0x5c7c32ed8730;  1 drivers
S_0x5c7c32ed6570 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ed6390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ed8730 .functor NAND 1, L_0x5c7c33122c40, L_0x5c7c33122ed0, C4<1>, C4<1>;
v0x5c7c32ed67c0_0 .net "in_a", 0 0, L_0x5c7c33122c40;  alias, 1 drivers
v0x5c7c32ed68a0_0 .net "in_b", 0 0, L_0x5c7c33122ed0;  alias, 1 drivers
v0x5c7c32ed6960_0 .net "out", 0 0, L_0x5c7c32ed8730;  alias, 1 drivers
S_0x5c7c32ed6ab0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ed6390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed7220_0 .net "in_a", 0 0, L_0x5c7c32ed8730;  alias, 1 drivers
v0x5c7c32ed72c0_0 .net "out", 0 0, L_0x5c7c331230b0;  alias, 1 drivers
S_0x5c7c32ed6cd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed6ab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331230b0 .functor NAND 1, L_0x5c7c32ed8730, L_0x5c7c32ed8730, C4<1>, C4<1>;
v0x5c7c32ed6f40_0 .net "in_a", 0 0, L_0x5c7c32ed8730;  alias, 1 drivers
v0x5c7c32ed7030_0 .net "in_b", 0 0, L_0x5c7c32ed8730;  alias, 1 drivers
v0x5c7c32ed7120_0 .net "out", 0 0, L_0x5c7c331230b0;  alias, 1 drivers
S_0x5c7c32ed77e0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32ed3950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed7f10_0 .net "in_a", 0 0, L_0x5c7c33122b90;  alias, 1 drivers
v0x5c7c32ed7fb0_0 .net "out", 0 0, L_0x5c7c33122c40;  alias, 1 drivers
S_0x5c7c32ed79b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed77e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122c40 .functor NAND 1, L_0x5c7c33122b90, L_0x5c7c33122b90, C4<1>, C4<1>;
v0x5c7c32ed7c20_0 .net "in_a", 0 0, L_0x5c7c33122b90;  alias, 1 drivers
v0x5c7c32ed7ce0_0 .net "in_b", 0 0, L_0x5c7c33122b90;  alias, 1 drivers
v0x5c7c32ed7e30_0 .net "out", 0 0, L_0x5c7c33122c40;  alias, 1 drivers
S_0x5c7c32ed80b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32ed3950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed8880_0 .net "in_a", 0 0, L_0x5c7c33122e20;  alias, 1 drivers
v0x5c7c32ed8920_0 .net "out", 0 0, L_0x5c7c33122ed0;  alias, 1 drivers
S_0x5c7c32ed8320 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed80b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33122ed0 .functor NAND 1, L_0x5c7c33122e20, L_0x5c7c33122e20, C4<1>, C4<1>;
v0x5c7c32ed8590_0 .net "in_a", 0 0, L_0x5c7c33122e20;  alias, 1 drivers
v0x5c7c32ed8650_0 .net "in_b", 0 0, L_0x5c7c33122e20;  alias, 1 drivers
v0x5c7c32ed87a0_0 .net "out", 0 0, L_0x5c7c33122ed0;  alias, 1 drivers
S_0x5c7c32ed8a20 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32ed3950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ed91c0_0 .net "in_a", 0 0, L_0x5c7c331230b0;  alias, 1 drivers
v0x5c7c32ed9260_0 .net "out", 0 0, L_0x5c7c33123160;  alias, 1 drivers
S_0x5c7c32ed8c40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ed8a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123160 .functor NAND 1, L_0x5c7c331230b0, L_0x5c7c331230b0, C4<1>, C4<1>;
v0x5c7c32ed8eb0_0 .net "in_a", 0 0, L_0x5c7c331230b0;  alias, 1 drivers
v0x5c7c32ed8f70_0 .net "in_b", 0 0, L_0x5c7c331230b0;  alias, 1 drivers
v0x5c7c32ed90c0_0 .net "out", 0 0, L_0x5c7c33123160;  alias, 1 drivers
S_0x5c7c32eda190 .scope module, "fa_gate9" "FullAdder" 2 14, 3 2 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /INPUT 1 "c";
    .port_info 3 /OUTPUT 1 "sum";
    .port_info 4 /OUTPUT 1 "carry";
v0x5c7c32ef8590_0 .net "a", 0 0, L_0x5c7c331259f0;  1 drivers
v0x5c7c32ef8630_0 .net "b", 0 0, L_0x5c7c33125a90;  1 drivers
v0x5c7c32ef86f0_0 .net "c", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ef8790_0 .net "carry", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32ef8830_0 .net "sum", 0 0, L_0x5c7c331250a0;  1 drivers
v0x5c7c32ef88d0_0 .net "tmp_carry_out_1", 0 0, L_0x5c7c33123660;  1 drivers
v0x5c7c32ef8970_0 .net "tmp_carry_out_2", 0 0, L_0x5c7c33124770;  1 drivers
v0x5c7c32ef8a10_0 .net "tmp_sum_out", 0 0, L_0x5c7c33124170;  1 drivers
S_0x5c7c32eda3f0 .scope module, "ha_gate1" "HalfAdder" 3 7, 4 3 0, S_0x5c7c32eda190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32ee5f70_0 .net "a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32ee6120_0 .net "b", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32ee62f0_0 .net "carry", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32ee6390_0 .net "sum", 0 0, L_0x5c7c33124170;  alias, 1 drivers
S_0x5c7c32eda660 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32eda3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32edb750_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edb820_0 .net "in_b", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32edb8f0_0 .net "out", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32edba10_0 .net "temp_out", 0 0, L_0x5c7c32ed9050;  1 drivers
S_0x5c7c32eda8d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32eda660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ed9050 .functor NAND 1, L_0x5c7c331259f0, L_0x5c7c33125a90, C4<1>, C4<1>;
v0x5c7c32edab40_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edac20_0 .net "in_b", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32edace0_0 .net "out", 0 0, L_0x5c7c32ed9050;  alias, 1 drivers
S_0x5c7c32edae30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32eda660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32edb5a0_0 .net "in_a", 0 0, L_0x5c7c32ed9050;  alias, 1 drivers
v0x5c7c32edb640_0 .net "out", 0 0, L_0x5c7c33123660;  alias, 1 drivers
S_0x5c7c32edb050 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32edae30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123660 .functor NAND 1, L_0x5c7c32ed9050, L_0x5c7c32ed9050, C4<1>, C4<1>;
v0x5c7c32edb2c0_0 .net "in_a", 0 0, L_0x5c7c32ed9050;  alias, 1 drivers
v0x5c7c32edb3b0_0 .net "in_b", 0 0, L_0x5c7c32ed9050;  alias, 1 drivers
v0x5c7c32edb4a0_0 .net "out", 0 0, L_0x5c7c33123660;  alias, 1 drivers
S_0x5c7c32edbad0 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32eda3f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee5890_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32ee5930_0 .net "in_b", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32ee59f0_0 .net "out", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ee5a90_0 .net "temp_a_and_out", 0 0, L_0x5c7c33123830;  1 drivers
v0x5c7c32ee5c40_0 .net "temp_a_out", 0 0, L_0x5c7c331236d0;  1 drivers
v0x5c7c32ee5ce0_0 .net "temp_b_and_out", 0 0, L_0x5c7c33123a40;  1 drivers
v0x5c7c32ee5e90_0 .net "temp_b_out", 0 0, L_0x5c7c331238e0;  1 drivers
S_0x5c7c32edbcb0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32edbad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32edcd70_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edce10_0 .net "in_b", 0 0, L_0x5c7c331236d0;  alias, 1 drivers
v0x5c7c32edcf00_0 .net "out", 0 0, L_0x5c7c33123830;  alias, 1 drivers
v0x5c7c32edd020_0 .net "temp_out", 0 0, L_0x5c7c33123780;  1 drivers
S_0x5c7c32edbf20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32edbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123780 .functor NAND 1, L_0x5c7c331259f0, L_0x5c7c331236d0, C4<1>, C4<1>;
v0x5c7c32edc190_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edc2a0_0 .net "in_b", 0 0, L_0x5c7c331236d0;  alias, 1 drivers
v0x5c7c32edc360_0 .net "out", 0 0, L_0x5c7c33123780;  alias, 1 drivers
S_0x5c7c32edc480 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32edbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32edcbc0_0 .net "in_a", 0 0, L_0x5c7c33123780;  alias, 1 drivers
v0x5c7c32edcc60_0 .net "out", 0 0, L_0x5c7c33123830;  alias, 1 drivers
S_0x5c7c32edc6a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32edc480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123830 .functor NAND 1, L_0x5c7c33123780, L_0x5c7c33123780, C4<1>, C4<1>;
v0x5c7c32edc910_0 .net "in_a", 0 0, L_0x5c7c33123780;  alias, 1 drivers
v0x5c7c32edc9d0_0 .net "in_b", 0 0, L_0x5c7c33123780;  alias, 1 drivers
v0x5c7c32edcac0_0 .net "out", 0 0, L_0x5c7c33123830;  alias, 1 drivers
S_0x5c7c32edd0e0 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32edbad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ede110_0 .net "in_a", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32ede1b0_0 .net "in_b", 0 0, L_0x5c7c331238e0;  alias, 1 drivers
v0x5c7c32ede2a0_0 .net "out", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
v0x5c7c32ede3c0_0 .net "temp_out", 0 0, L_0x5c7c33123990;  1 drivers
S_0x5c7c32edd2c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32edd0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123990 .functor NAND 1, L_0x5c7c33125a90, L_0x5c7c331238e0, C4<1>, C4<1>;
v0x5c7c32edd530_0 .net "in_a", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32edd640_0 .net "in_b", 0 0, L_0x5c7c331238e0;  alias, 1 drivers
v0x5c7c32edd700_0 .net "out", 0 0, L_0x5c7c33123990;  alias, 1 drivers
S_0x5c7c32edd820 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32edd0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eddf60_0 .net "in_a", 0 0, L_0x5c7c33123990;  alias, 1 drivers
v0x5c7c32ede000_0 .net "out", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
S_0x5c7c32edda40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32edd820;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123a40 .functor NAND 1, L_0x5c7c33123990, L_0x5c7c33123990, C4<1>, C4<1>;
v0x5c7c32eddcb0_0 .net "in_a", 0 0, L_0x5c7c33123990;  alias, 1 drivers
v0x5c7c32eddd70_0 .net "in_b", 0 0, L_0x5c7c33123990;  alias, 1 drivers
v0x5c7c32edde60_0 .net "out", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
S_0x5c7c32ede510 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32edbad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32edec50_0 .net "in_a", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32edecf0_0 .net "out", 0 0, L_0x5c7c331236d0;  alias, 1 drivers
S_0x5c7c32ede6e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ede510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331236d0 .functor NAND 1, L_0x5c7c33125a90, L_0x5c7c33125a90, C4<1>, C4<1>;
v0x5c7c32ede930_0 .net "in_a", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32edea80_0 .net "in_b", 0 0, L_0x5c7c33125a90;  alias, 1 drivers
v0x5c7c32edeb40_0 .net "out", 0 0, L_0x5c7c331236d0;  alias, 1 drivers
S_0x5c7c32ededf0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32edbad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32edf570_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edf610_0 .net "out", 0 0, L_0x5c7c331238e0;  alias, 1 drivers
S_0x5c7c32edf010 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ededf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331238e0 .functor NAND 1, L_0x5c7c331259f0, L_0x5c7c331259f0, C4<1>, C4<1>;
v0x5c7c32edf280_0 .net "in_a", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edf3d0_0 .net "in_b", 0 0, L_0x5c7c331259f0;  alias, 1 drivers
v0x5c7c32edf490_0 .net "out", 0 0, L_0x5c7c331238e0;  alias, 1 drivers
S_0x5c7c32edf710 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32edbad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee51e0_0 .net "branch1_out", 0 0, L_0x5c7c33123c50;  1 drivers
v0x5c7c32ee5310_0 .net "branch2_out", 0 0, L_0x5c7c33123ee0;  1 drivers
v0x5c7c32ee5460_0 .net "in_a", 0 0, L_0x5c7c33123830;  alias, 1 drivers
v0x5c7c32ee5530_0 .net "in_b", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
v0x5c7c32ee55d0_0 .net "out", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ee5670_0 .net "temp1_out", 0 0, L_0x5c7c33123ba0;  1 drivers
v0x5c7c32ee5710_0 .net "temp2_out", 0 0, L_0x5c7c33123e30;  1 drivers
v0x5c7c32ee57b0_0 .net "temp3_out", 0 0, L_0x5c7c331240c0;  1 drivers
S_0x5c7c32edf990 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32edf710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee0a20_0 .net "in_a", 0 0, L_0x5c7c33123830;  alias, 1 drivers
v0x5c7c32ee0ac0_0 .net "in_b", 0 0, L_0x5c7c33123830;  alias, 1 drivers
v0x5c7c32ee0b80_0 .net "out", 0 0, L_0x5c7c33123ba0;  alias, 1 drivers
v0x5c7c32ee0ca0_0 .net "temp_out", 0 0, L_0x5c7c33123af0;  1 drivers
S_0x5c7c32edfc00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32edf990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123af0 .functor NAND 1, L_0x5c7c33123830, L_0x5c7c33123830, C4<1>, C4<1>;
v0x5c7c32edfe70_0 .net "in_a", 0 0, L_0x5c7c33123830;  alias, 1 drivers
v0x5c7c32edff30_0 .net "in_b", 0 0, L_0x5c7c33123830;  alias, 1 drivers
v0x5c7c32ee0080_0 .net "out", 0 0, L_0x5c7c33123af0;  alias, 1 drivers
S_0x5c7c32ee0180 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32edf990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee0870_0 .net "in_a", 0 0, L_0x5c7c33123af0;  alias, 1 drivers
v0x5c7c32ee0910_0 .net "out", 0 0, L_0x5c7c33123ba0;  alias, 1 drivers
S_0x5c7c32ee0350 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee0180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123ba0 .functor NAND 1, L_0x5c7c33123af0, L_0x5c7c33123af0, C4<1>, C4<1>;
v0x5c7c32ee05c0_0 .net "in_a", 0 0, L_0x5c7c33123af0;  alias, 1 drivers
v0x5c7c32ee0680_0 .net "in_b", 0 0, L_0x5c7c33123af0;  alias, 1 drivers
v0x5c7c32ee0770_0 .net "out", 0 0, L_0x5c7c33123ba0;  alias, 1 drivers
S_0x5c7c32ee0e10 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32edf710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee1e40_0 .net "in_a", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
v0x5c7c32ee1ee0_0 .net "in_b", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
v0x5c7c32ee1fa0_0 .net "out", 0 0, L_0x5c7c33123e30;  alias, 1 drivers
v0x5c7c32ee20c0_0 .net "temp_out", 0 0, L_0x5c7c32ee3c60;  1 drivers
S_0x5c7c32ee0ff0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ee0e10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ee3c60 .functor NAND 1, L_0x5c7c33123a40, L_0x5c7c33123a40, C4<1>, C4<1>;
v0x5c7c32ee1260_0 .net "in_a", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
v0x5c7c32ee1320_0 .net "in_b", 0 0, L_0x5c7c33123a40;  alias, 1 drivers
v0x5c7c32ee1470_0 .net "out", 0 0, L_0x5c7c32ee3c60;  alias, 1 drivers
S_0x5c7c32ee1570 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ee0e10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee1c90_0 .net "in_a", 0 0, L_0x5c7c32ee3c60;  alias, 1 drivers
v0x5c7c32ee1d30_0 .net "out", 0 0, L_0x5c7c33123e30;  alias, 1 drivers
S_0x5c7c32ee1740 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee1570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123e30 .functor NAND 1, L_0x5c7c32ee3c60, L_0x5c7c32ee3c60, C4<1>, C4<1>;
v0x5c7c32ee19b0_0 .net "in_a", 0 0, L_0x5c7c32ee3c60;  alias, 1 drivers
v0x5c7c32ee1aa0_0 .net "in_b", 0 0, L_0x5c7c32ee3c60;  alias, 1 drivers
v0x5c7c32ee1b90_0 .net "out", 0 0, L_0x5c7c33123e30;  alias, 1 drivers
S_0x5c7c32ee2230 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32edf710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee3270_0 .net "in_a", 0 0, L_0x5c7c33123c50;  alias, 1 drivers
v0x5c7c32ee3340_0 .net "in_b", 0 0, L_0x5c7c33123ee0;  alias, 1 drivers
v0x5c7c32ee3410_0 .net "out", 0 0, L_0x5c7c331240c0;  alias, 1 drivers
v0x5c7c32ee3530_0 .net "temp_out", 0 0, L_0x5c7c32ee45d0;  1 drivers
S_0x5c7c32ee2410 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ee2230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ee45d0 .functor NAND 1, L_0x5c7c33123c50, L_0x5c7c33123ee0, C4<1>, C4<1>;
v0x5c7c32ee2660_0 .net "in_a", 0 0, L_0x5c7c33123c50;  alias, 1 drivers
v0x5c7c32ee2740_0 .net "in_b", 0 0, L_0x5c7c33123ee0;  alias, 1 drivers
v0x5c7c32ee2800_0 .net "out", 0 0, L_0x5c7c32ee45d0;  alias, 1 drivers
S_0x5c7c32ee2950 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ee2230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee30c0_0 .net "in_a", 0 0, L_0x5c7c32ee45d0;  alias, 1 drivers
v0x5c7c32ee3160_0 .net "out", 0 0, L_0x5c7c331240c0;  alias, 1 drivers
S_0x5c7c32ee2b70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee2950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331240c0 .functor NAND 1, L_0x5c7c32ee45d0, L_0x5c7c32ee45d0, C4<1>, C4<1>;
v0x5c7c32ee2de0_0 .net "in_a", 0 0, L_0x5c7c32ee45d0;  alias, 1 drivers
v0x5c7c32ee2ed0_0 .net "in_b", 0 0, L_0x5c7c32ee45d0;  alias, 1 drivers
v0x5c7c32ee2fc0_0 .net "out", 0 0, L_0x5c7c331240c0;  alias, 1 drivers
S_0x5c7c32ee3680 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32edf710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee3db0_0 .net "in_a", 0 0, L_0x5c7c33123ba0;  alias, 1 drivers
v0x5c7c32ee3e50_0 .net "out", 0 0, L_0x5c7c33123c50;  alias, 1 drivers
S_0x5c7c32ee3850 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee3680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123c50 .functor NAND 1, L_0x5c7c33123ba0, L_0x5c7c33123ba0, C4<1>, C4<1>;
v0x5c7c32ee3ac0_0 .net "in_a", 0 0, L_0x5c7c33123ba0;  alias, 1 drivers
v0x5c7c32ee3b80_0 .net "in_b", 0 0, L_0x5c7c33123ba0;  alias, 1 drivers
v0x5c7c32ee3cd0_0 .net "out", 0 0, L_0x5c7c33123c50;  alias, 1 drivers
S_0x5c7c32ee3f50 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32edf710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee4720_0 .net "in_a", 0 0, L_0x5c7c33123e30;  alias, 1 drivers
v0x5c7c32ee47c0_0 .net "out", 0 0, L_0x5c7c33123ee0;  alias, 1 drivers
S_0x5c7c32ee41c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee3f50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33123ee0 .functor NAND 1, L_0x5c7c33123e30, L_0x5c7c33123e30, C4<1>, C4<1>;
v0x5c7c32ee4430_0 .net "in_a", 0 0, L_0x5c7c33123e30;  alias, 1 drivers
v0x5c7c32ee44f0_0 .net "in_b", 0 0, L_0x5c7c33123e30;  alias, 1 drivers
v0x5c7c32ee4640_0 .net "out", 0 0, L_0x5c7c33123ee0;  alias, 1 drivers
S_0x5c7c32ee48c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32edf710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee5060_0 .net "in_a", 0 0, L_0x5c7c331240c0;  alias, 1 drivers
v0x5c7c32ee5100_0 .net "out", 0 0, L_0x5c7c33124170;  alias, 1 drivers
S_0x5c7c32ee4ae0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee48c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124170 .functor NAND 1, L_0x5c7c331240c0, L_0x5c7c331240c0, C4<1>, C4<1>;
v0x5c7c32ee4d50_0 .net "in_a", 0 0, L_0x5c7c331240c0;  alias, 1 drivers
v0x5c7c32ee4e10_0 .net "in_b", 0 0, L_0x5c7c331240c0;  alias, 1 drivers
v0x5c7c32ee4f60_0 .net "out", 0 0, L_0x5c7c33124170;  alias, 1 drivers
S_0x5c7c32ee6470 .scope module, "ha_gate2" "HalfAdder" 3 8, 4 3 0, S_0x5c7c32eda190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32ef1f90_0 .net "a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ef2030_0 .net "b", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ef20f0_0 .net "carry", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ef2190_0 .net "sum", 0 0, L_0x5c7c331250a0;  alias, 1 drivers
S_0x5c7c32ee6690 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32ee6470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee7630_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ee76d0_0 .net "in_b", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ee7790_0 .net "out", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ee78b0_0 .net "temp_out", 0 0, L_0x5c7c32ee4ef0;  1 drivers
S_0x5c7c32ee6840 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ee6690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ee4ef0 .functor NAND 1, L_0x5c7c33124170, L_0x5c7c33123160, C4<1>, C4<1>;
v0x5c7c32ee6ab0_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ee6b70_0 .net "in_b", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ee6c30_0 .net "out", 0 0, L_0x5c7c32ee4ef0;  alias, 1 drivers
S_0x5c7c32ee6d60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ee6690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee7480_0 .net "in_a", 0 0, L_0x5c7c32ee4ef0;  alias, 1 drivers
v0x5c7c32ee7520_0 .net "out", 0 0, L_0x5c7c33124770;  alias, 1 drivers
S_0x5c7c32ee6f30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee6d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124770 .functor NAND 1, L_0x5c7c32ee4ef0, L_0x5c7c32ee4ef0, C4<1>, C4<1>;
v0x5c7c32ee71a0_0 .net "in_a", 0 0, L_0x5c7c32ee4ef0;  alias, 1 drivers
v0x5c7c32ee7290_0 .net "in_b", 0 0, L_0x5c7c32ee4ef0;  alias, 1 drivers
v0x5c7c32ee7380_0 .net "out", 0 0, L_0x5c7c33124770;  alias, 1 drivers
S_0x5c7c32ee7a20 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32ee6470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef18b0_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ef1950_0 .net "in_b", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ef1a10_0 .net "out", 0 0, L_0x5c7c331250a0;  alias, 1 drivers
v0x5c7c32ef1ab0_0 .net "temp_a_and_out", 0 0, L_0x5c7c33124980;  1 drivers
v0x5c7c32ef1c60_0 .net "temp_a_out", 0 0, L_0x5c7c33124820;  1 drivers
v0x5c7c32ef1d00_0 .net "temp_b_and_out", 0 0, L_0x5c7c33124b90;  1 drivers
v0x5c7c32ef1eb0_0 .net "temp_b_out", 0 0, L_0x5c7c33124a30;  1 drivers
S_0x5c7c32ee7c00 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32ee7a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ee8ca0_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ee8e50_0 .net "in_b", 0 0, L_0x5c7c33124820;  alias, 1 drivers
v0x5c7c32ee8f40_0 .net "out", 0 0, L_0x5c7c33124980;  alias, 1 drivers
v0x5c7c32ee9060_0 .net "temp_out", 0 0, L_0x5c7c331248d0;  1 drivers
S_0x5c7c32ee7e70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ee7c00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331248d0 .functor NAND 1, L_0x5c7c33124170, L_0x5c7c33124820, C4<1>, C4<1>;
v0x5c7c32ee80e0_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32ee81a0_0 .net "in_b", 0 0, L_0x5c7c33124820;  alias, 1 drivers
v0x5c7c32ee8260_0 .net "out", 0 0, L_0x5c7c331248d0;  alias, 1 drivers
S_0x5c7c32ee8380 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ee7c00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee8af0_0 .net "in_a", 0 0, L_0x5c7c331248d0;  alias, 1 drivers
v0x5c7c32ee8b90_0 .net "out", 0 0, L_0x5c7c33124980;  alias, 1 drivers
S_0x5c7c32ee85a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee8380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124980 .functor NAND 1, L_0x5c7c331248d0, L_0x5c7c331248d0, C4<1>, C4<1>;
v0x5c7c32ee8810_0 .net "in_a", 0 0, L_0x5c7c331248d0;  alias, 1 drivers
v0x5c7c32ee8900_0 .net "in_b", 0 0, L_0x5c7c331248d0;  alias, 1 drivers
v0x5c7c32ee89f0_0 .net "out", 0 0, L_0x5c7c33124980;  alias, 1 drivers
S_0x5c7c32ee9120 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32ee7a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32eea130_0 .net "in_a", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32eea1d0_0 .net "in_b", 0 0, L_0x5c7c33124a30;  alias, 1 drivers
v0x5c7c32eea2c0_0 .net "out", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
v0x5c7c32eea3e0_0 .net "temp_out", 0 0, L_0x5c7c33124ae0;  1 drivers
S_0x5c7c32ee9300 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ee9120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124ae0 .functor NAND 1, L_0x5c7c33123160, L_0x5c7c33124a30, C4<1>, C4<1>;
v0x5c7c32ee9570_0 .net "in_a", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32ee9630_0 .net "in_b", 0 0, L_0x5c7c33124a30;  alias, 1 drivers
v0x5c7c32ee96f0_0 .net "out", 0 0, L_0x5c7c33124ae0;  alias, 1 drivers
S_0x5c7c32ee9810 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ee9120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ee9f80_0 .net "in_a", 0 0, L_0x5c7c33124ae0;  alias, 1 drivers
v0x5c7c32eea020_0 .net "out", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
S_0x5c7c32ee9a30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ee9810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124b90 .functor NAND 1, L_0x5c7c33124ae0, L_0x5c7c33124ae0, C4<1>, C4<1>;
v0x5c7c32ee9ca0_0 .net "in_a", 0 0, L_0x5c7c33124ae0;  alias, 1 drivers
v0x5c7c32ee9d90_0 .net "in_b", 0 0, L_0x5c7c33124ae0;  alias, 1 drivers
v0x5c7c32ee9e80_0 .net "out", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
S_0x5c7c32eea530 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32ee7a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eead40_0 .net "in_a", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32eeade0_0 .net "out", 0 0, L_0x5c7c33124820;  alias, 1 drivers
S_0x5c7c32eea700 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eea530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124820 .functor NAND 1, L_0x5c7c33123160, L_0x5c7c33123160, C4<1>, C4<1>;
v0x5c7c32eea950_0 .net "in_a", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32eeab20_0 .net "in_b", 0 0, L_0x5c7c33123160;  alias, 1 drivers
v0x5c7c32eeabe0_0 .net "out", 0 0, L_0x5c7c33124820;  alias, 1 drivers
S_0x5c7c32eeaee0 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32ee7a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eeb620_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32eeb6c0_0 .net "out", 0 0, L_0x5c7c33124a30;  alias, 1 drivers
S_0x5c7c32eeb100 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eeaee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124a30 .functor NAND 1, L_0x5c7c33124170, L_0x5c7c33124170, C4<1>, C4<1>;
v0x5c7c32eeb370_0 .net "in_a", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32eeb430_0 .net "in_b", 0 0, L_0x5c7c33124170;  alias, 1 drivers
v0x5c7c32eeb4f0_0 .net "out", 0 0, L_0x5c7c33124a30;  alias, 1 drivers
S_0x5c7c32eeb7c0 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32ee7a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef1200_0 .net "branch1_out", 0 0, L_0x5c7c33124da0;  1 drivers
v0x5c7c32ef1330_0 .net "branch2_out", 0 0, L_0x5c7c33124f20;  1 drivers
v0x5c7c32ef1480_0 .net "in_a", 0 0, L_0x5c7c33124980;  alias, 1 drivers
v0x5c7c32ef1550_0 .net "in_b", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
v0x5c7c32ef15f0_0 .net "out", 0 0, L_0x5c7c331250a0;  alias, 1 drivers
v0x5c7c32ef1690_0 .net "temp1_out", 0 0, L_0x5c7c33124cf0;  1 drivers
v0x5c7c32ef1730_0 .net "temp2_out", 0 0, L_0x5c7c33124e70;  1 drivers
v0x5c7c32ef17d0_0 .net "temp3_out", 0 0, L_0x5c7c33124ff0;  1 drivers
S_0x5c7c32eeba40 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32eeb7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32eeca40_0 .net "in_a", 0 0, L_0x5c7c33124980;  alias, 1 drivers
v0x5c7c32eecae0_0 .net "in_b", 0 0, L_0x5c7c33124980;  alias, 1 drivers
v0x5c7c32eecba0_0 .net "out", 0 0, L_0x5c7c33124cf0;  alias, 1 drivers
v0x5c7c32eeccc0_0 .net "temp_out", 0 0, L_0x5c7c33124c40;  1 drivers
S_0x5c7c32eebcb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32eeba40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124c40 .functor NAND 1, L_0x5c7c33124980, L_0x5c7c33124980, C4<1>, C4<1>;
v0x5c7c32eebf20_0 .net "in_a", 0 0, L_0x5c7c33124980;  alias, 1 drivers
v0x5c7c32eebfe0_0 .net "in_b", 0 0, L_0x5c7c33124980;  alias, 1 drivers
v0x5c7c32eec0a0_0 .net "out", 0 0, L_0x5c7c33124c40;  alias, 1 drivers
S_0x5c7c32eec1a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32eeba40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eec890_0 .net "in_a", 0 0, L_0x5c7c33124c40;  alias, 1 drivers
v0x5c7c32eec930_0 .net "out", 0 0, L_0x5c7c33124cf0;  alias, 1 drivers
S_0x5c7c32eec370 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eec1a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124cf0 .functor NAND 1, L_0x5c7c33124c40, L_0x5c7c33124c40, C4<1>, C4<1>;
v0x5c7c32eec5e0_0 .net "in_a", 0 0, L_0x5c7c33124c40;  alias, 1 drivers
v0x5c7c32eec6a0_0 .net "in_b", 0 0, L_0x5c7c33124c40;  alias, 1 drivers
v0x5c7c32eec790_0 .net "out", 0 0, L_0x5c7c33124cf0;  alias, 1 drivers
S_0x5c7c32eece30 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32eeb7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32eede60_0 .net "in_a", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
v0x5c7c32eedf00_0 .net "in_b", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
v0x5c7c32eedfc0_0 .net "out", 0 0, L_0x5c7c33124e70;  alias, 1 drivers
v0x5c7c32eee0e0_0 .net "temp_out", 0 0, L_0x5c7c32eefc80;  1 drivers
S_0x5c7c32eed010 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32eece30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32eefc80 .functor NAND 1, L_0x5c7c33124b90, L_0x5c7c33124b90, C4<1>, C4<1>;
v0x5c7c32eed280_0 .net "in_a", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
v0x5c7c32eed340_0 .net "in_b", 0 0, L_0x5c7c33124b90;  alias, 1 drivers
v0x5c7c32eed490_0 .net "out", 0 0, L_0x5c7c32eefc80;  alias, 1 drivers
S_0x5c7c32eed590 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32eece30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eedcb0_0 .net "in_a", 0 0, L_0x5c7c32eefc80;  alias, 1 drivers
v0x5c7c32eedd50_0 .net "out", 0 0, L_0x5c7c33124e70;  alias, 1 drivers
S_0x5c7c32eed760 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eed590;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124e70 .functor NAND 1, L_0x5c7c32eefc80, L_0x5c7c32eefc80, C4<1>, C4<1>;
v0x5c7c32eed9d0_0 .net "in_a", 0 0, L_0x5c7c32eefc80;  alias, 1 drivers
v0x5c7c32eedac0_0 .net "in_b", 0 0, L_0x5c7c32eefc80;  alias, 1 drivers
v0x5c7c32eedbb0_0 .net "out", 0 0, L_0x5c7c33124e70;  alias, 1 drivers
S_0x5c7c32eee250 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32eeb7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32eef290_0 .net "in_a", 0 0, L_0x5c7c33124da0;  alias, 1 drivers
v0x5c7c32eef360_0 .net "in_b", 0 0, L_0x5c7c33124f20;  alias, 1 drivers
v0x5c7c32eef430_0 .net "out", 0 0, L_0x5c7c33124ff0;  alias, 1 drivers
v0x5c7c32eef550_0 .net "temp_out", 0 0, L_0x5c7c32ef05f0;  1 drivers
S_0x5c7c32eee430 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32eee250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ef05f0 .functor NAND 1, L_0x5c7c33124da0, L_0x5c7c33124f20, C4<1>, C4<1>;
v0x5c7c32eee680_0 .net "in_a", 0 0, L_0x5c7c33124da0;  alias, 1 drivers
v0x5c7c32eee760_0 .net "in_b", 0 0, L_0x5c7c33124f20;  alias, 1 drivers
v0x5c7c32eee820_0 .net "out", 0 0, L_0x5c7c32ef05f0;  alias, 1 drivers
S_0x5c7c32eee970 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32eee250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eef0e0_0 .net "in_a", 0 0, L_0x5c7c32ef05f0;  alias, 1 drivers
v0x5c7c32eef180_0 .net "out", 0 0, L_0x5c7c33124ff0;  alias, 1 drivers
S_0x5c7c32eeeb90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eee970;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124ff0 .functor NAND 1, L_0x5c7c32ef05f0, L_0x5c7c32ef05f0, C4<1>, C4<1>;
v0x5c7c32eeee00_0 .net "in_a", 0 0, L_0x5c7c32ef05f0;  alias, 1 drivers
v0x5c7c32eeeef0_0 .net "in_b", 0 0, L_0x5c7c32ef05f0;  alias, 1 drivers
v0x5c7c32eeefe0_0 .net "out", 0 0, L_0x5c7c33124ff0;  alias, 1 drivers
S_0x5c7c32eef6a0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32eeb7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32eefdd0_0 .net "in_a", 0 0, L_0x5c7c33124cf0;  alias, 1 drivers
v0x5c7c32eefe70_0 .net "out", 0 0, L_0x5c7c33124da0;  alias, 1 drivers
S_0x5c7c32eef870 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eef6a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124da0 .functor NAND 1, L_0x5c7c33124cf0, L_0x5c7c33124cf0, C4<1>, C4<1>;
v0x5c7c32eefae0_0 .net "in_a", 0 0, L_0x5c7c33124cf0;  alias, 1 drivers
v0x5c7c32eefba0_0 .net "in_b", 0 0, L_0x5c7c33124cf0;  alias, 1 drivers
v0x5c7c32eefcf0_0 .net "out", 0 0, L_0x5c7c33124da0;  alias, 1 drivers
S_0x5c7c32eeff70 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32eeb7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef0740_0 .net "in_a", 0 0, L_0x5c7c33124e70;  alias, 1 drivers
v0x5c7c32ef07e0_0 .net "out", 0 0, L_0x5c7c33124f20;  alias, 1 drivers
S_0x5c7c32ef01e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32eeff70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33124f20 .functor NAND 1, L_0x5c7c33124e70, L_0x5c7c33124e70, C4<1>, C4<1>;
v0x5c7c32ef0450_0 .net "in_a", 0 0, L_0x5c7c33124e70;  alias, 1 drivers
v0x5c7c32ef0510_0 .net "in_b", 0 0, L_0x5c7c33124e70;  alias, 1 drivers
v0x5c7c32ef0660_0 .net "out", 0 0, L_0x5c7c33124f20;  alias, 1 drivers
S_0x5c7c32ef08e0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32eeb7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef1080_0 .net "in_a", 0 0, L_0x5c7c33124ff0;  alias, 1 drivers
v0x5c7c32ef1120_0 .net "out", 0 0, L_0x5c7c331250a0;  alias, 1 drivers
S_0x5c7c32ef0b00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef08e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331250a0 .functor NAND 1, L_0x5c7c33124ff0, L_0x5c7c33124ff0, C4<1>, C4<1>;
v0x5c7c32ef0d70_0 .net "in_a", 0 0, L_0x5c7c33124ff0;  alias, 1 drivers
v0x5c7c32ef0e30_0 .net "in_b", 0 0, L_0x5c7c33124ff0;  alias, 1 drivers
v0x5c7c32ef0f80_0 .net "out", 0 0, L_0x5c7c331250a0;  alias, 1 drivers
S_0x5c7c32ef2300 .scope module, "or_gate" "Or" 3 9, 9 3 0, S_0x5c7c32eda190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef7cf0_0 .net "branch1_out", 0 0, L_0x5c7c33125330;  1 drivers
v0x5c7c32ef7e20_0 .net "branch2_out", 0 0, L_0x5c7c331255c0;  1 drivers
v0x5c7c32ef7f70_0 .net "in_a", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32ef8120_0 .net "in_b", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ef82d0_0 .net "out", 0 0, L_0x5c7c33125850;  alias, 1 drivers
v0x5c7c32ef8370_0 .net "temp1_out", 0 0, L_0x5c7c33125280;  1 drivers
v0x5c7c32ef8410_0 .net "temp2_out", 0 0, L_0x5c7c33125510;  1 drivers
v0x5c7c32ef84b0_0 .net "temp3_out", 0 0, L_0x5c7c331257a0;  1 drivers
S_0x5c7c32ef2490 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32ef2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef3530_0 .net "in_a", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32ef35d0_0 .net "in_b", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32ef3690_0 .net "out", 0 0, L_0x5c7c33125280;  alias, 1 drivers
v0x5c7c32ef37b0_0 .net "temp_out", 0 0, L_0x5c7c32ef0f10;  1 drivers
S_0x5c7c32ef26b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ef2490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ef0f10 .functor NAND 1, L_0x5c7c33123660, L_0x5c7c33123660, C4<1>, C4<1>;
v0x5c7c32ef2920_0 .net "in_a", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32ef2a70_0 .net "in_b", 0 0, L_0x5c7c33123660;  alias, 1 drivers
v0x5c7c32ef2b30_0 .net "out", 0 0, L_0x5c7c32ef0f10;  alias, 1 drivers
S_0x5c7c32ef2c60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ef2490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef3380_0 .net "in_a", 0 0, L_0x5c7c32ef0f10;  alias, 1 drivers
v0x5c7c32ef3420_0 .net "out", 0 0, L_0x5c7c33125280;  alias, 1 drivers
S_0x5c7c32ef2e30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef2c60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125280 .functor NAND 1, L_0x5c7c32ef0f10, L_0x5c7c32ef0f10, C4<1>, C4<1>;
v0x5c7c32ef30a0_0 .net "in_a", 0 0, L_0x5c7c32ef0f10;  alias, 1 drivers
v0x5c7c32ef3190_0 .net "in_b", 0 0, L_0x5c7c32ef0f10;  alias, 1 drivers
v0x5c7c32ef3280_0 .net "out", 0 0, L_0x5c7c33125280;  alias, 1 drivers
S_0x5c7c32ef3920 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32ef2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef4950_0 .net "in_a", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ef49f0_0 .net "in_b", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ef4ab0_0 .net "out", 0 0, L_0x5c7c33125510;  alias, 1 drivers
v0x5c7c32ef4bd0_0 .net "temp_out", 0 0, L_0x5c7c32ef6770;  1 drivers
S_0x5c7c32ef3b00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ef3920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ef6770 .functor NAND 1, L_0x5c7c33124770, L_0x5c7c33124770, C4<1>, C4<1>;
v0x5c7c32ef3d70_0 .net "in_a", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ef3ec0_0 .net "in_b", 0 0, L_0x5c7c33124770;  alias, 1 drivers
v0x5c7c32ef3f80_0 .net "out", 0 0, L_0x5c7c32ef6770;  alias, 1 drivers
S_0x5c7c32ef4080 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ef3920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef47a0_0 .net "in_a", 0 0, L_0x5c7c32ef6770;  alias, 1 drivers
v0x5c7c32ef4840_0 .net "out", 0 0, L_0x5c7c33125510;  alias, 1 drivers
S_0x5c7c32ef4250 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef4080;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125510 .functor NAND 1, L_0x5c7c32ef6770, L_0x5c7c32ef6770, C4<1>, C4<1>;
v0x5c7c32ef44c0_0 .net "in_a", 0 0, L_0x5c7c32ef6770;  alias, 1 drivers
v0x5c7c32ef45b0_0 .net "in_b", 0 0, L_0x5c7c32ef6770;  alias, 1 drivers
v0x5c7c32ef46a0_0 .net "out", 0 0, L_0x5c7c33125510;  alias, 1 drivers
S_0x5c7c32ef4d40 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32ef2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef5d80_0 .net "in_a", 0 0, L_0x5c7c33125330;  alias, 1 drivers
v0x5c7c32ef5e50_0 .net "in_b", 0 0, L_0x5c7c331255c0;  alias, 1 drivers
v0x5c7c32ef5f20_0 .net "out", 0 0, L_0x5c7c331257a0;  alias, 1 drivers
v0x5c7c32ef6040_0 .net "temp_out", 0 0, L_0x5c7c32ef70e0;  1 drivers
S_0x5c7c32ef4f20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ef4d40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32ef70e0 .functor NAND 1, L_0x5c7c33125330, L_0x5c7c331255c0, C4<1>, C4<1>;
v0x5c7c32ef5170_0 .net "in_a", 0 0, L_0x5c7c33125330;  alias, 1 drivers
v0x5c7c32ef5250_0 .net "in_b", 0 0, L_0x5c7c331255c0;  alias, 1 drivers
v0x5c7c32ef5310_0 .net "out", 0 0, L_0x5c7c32ef70e0;  alias, 1 drivers
S_0x5c7c32ef5460 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ef4d40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef5bd0_0 .net "in_a", 0 0, L_0x5c7c32ef70e0;  alias, 1 drivers
v0x5c7c32ef5c70_0 .net "out", 0 0, L_0x5c7c331257a0;  alias, 1 drivers
S_0x5c7c32ef5680 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef5460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331257a0 .functor NAND 1, L_0x5c7c32ef70e0, L_0x5c7c32ef70e0, C4<1>, C4<1>;
v0x5c7c32ef58f0_0 .net "in_a", 0 0, L_0x5c7c32ef70e0;  alias, 1 drivers
v0x5c7c32ef59e0_0 .net "in_b", 0 0, L_0x5c7c32ef70e0;  alias, 1 drivers
v0x5c7c32ef5ad0_0 .net "out", 0 0, L_0x5c7c331257a0;  alias, 1 drivers
S_0x5c7c32ef6190 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32ef2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef68c0_0 .net "in_a", 0 0, L_0x5c7c33125280;  alias, 1 drivers
v0x5c7c32ef6960_0 .net "out", 0 0, L_0x5c7c33125330;  alias, 1 drivers
S_0x5c7c32ef6360 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef6190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125330 .functor NAND 1, L_0x5c7c33125280, L_0x5c7c33125280, C4<1>, C4<1>;
v0x5c7c32ef65d0_0 .net "in_a", 0 0, L_0x5c7c33125280;  alias, 1 drivers
v0x5c7c32ef6690_0 .net "in_b", 0 0, L_0x5c7c33125280;  alias, 1 drivers
v0x5c7c32ef67e0_0 .net "out", 0 0, L_0x5c7c33125330;  alias, 1 drivers
S_0x5c7c32ef6a60 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32ef2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef7230_0 .net "in_a", 0 0, L_0x5c7c33125510;  alias, 1 drivers
v0x5c7c32ef72d0_0 .net "out", 0 0, L_0x5c7c331255c0;  alias, 1 drivers
S_0x5c7c32ef6cd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef6a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331255c0 .functor NAND 1, L_0x5c7c33125510, L_0x5c7c33125510, C4<1>, C4<1>;
v0x5c7c32ef6f40_0 .net "in_a", 0 0, L_0x5c7c33125510;  alias, 1 drivers
v0x5c7c32ef7000_0 .net "in_b", 0 0, L_0x5c7c33125510;  alias, 1 drivers
v0x5c7c32ef7150_0 .net "out", 0 0, L_0x5c7c331255c0;  alias, 1 drivers
S_0x5c7c32ef73d0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32ef2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef7b50_0 .net "in_a", 0 0, L_0x5c7c331257a0;  alias, 1 drivers
v0x5c7c32ef7bf0_0 .net "out", 0 0, L_0x5c7c33125850;  alias, 1 drivers
S_0x5c7c32ef75f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef73d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33125850 .functor NAND 1, L_0x5c7c331257a0, L_0x5c7c331257a0, C4<1>, C4<1>;
v0x5c7c32ef7860_0 .net "in_a", 0 0, L_0x5c7c331257a0;  alias, 1 drivers
v0x5c7c32ef7920_0 .net "in_b", 0 0, L_0x5c7c331257a0;  alias, 1 drivers
v0x5c7c32ef7a70_0 .net "out", 0 0, L_0x5c7c33125850;  alias, 1 drivers
S_0x5c7c32ef8b10 .scope module, "ha_gate1" "HalfAdder" 2 6, 4 3 0, S_0x5c7c329f9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "a";
    .port_info 1 /INPUT 1 "b";
    .port_info 2 /OUTPUT 1 "sum";
    .port_info 3 /OUTPUT 1 "carry";
v0x5c7c32f045d0_0 .net "a", 0 0, L_0x5c7c33112b10;  1 drivers
v0x5c7c32f04780_0 .net "b", 0 0, L_0x5c7c33112be0;  1 drivers
v0x5c7c32f04950_0 .net "carry", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32f049f0_0 .net "sum", 0 0, L_0x5c7c33112950;  1 drivers
S_0x5c7c32ef8d10 .scope module, "and_gate" "And" 4 7, 5 2 0, S_0x5c7c32ef8b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ef9dd0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32ef9ea0_0 .net "in_b", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32ef9f70_0 .net "out", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
v0x5c7c32efa040_0 .net "temp_out", 0 0, L_0x5c7c33111c30;  1 drivers
S_0x5c7c32ef8f80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ef8d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33111c30 .functor NAND 1, L_0x5c7c33112b10, L_0x5c7c33112be0, C4<1>, C4<1>;
v0x5c7c32ef91f0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32ef92d0_0 .net "in_b", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32ef9390_0 .net "out", 0 0, L_0x5c7c33111c30;  alias, 1 drivers
S_0x5c7c32ef94e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ef8d10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ef9c30_0 .net "in_a", 0 0, L_0x5c7c33111c30;  alias, 1 drivers
v0x5c7c32ef9cd0_0 .net "out", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
S_0x5c7c32ef9700 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ef94e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33111ce0 .functor NAND 1, L_0x5c7c33111c30, L_0x5c7c33111c30, C4<1>, C4<1>;
v0x5c7c32ef9970_0 .net "in_a", 0 0, L_0x5c7c33111c30;  alias, 1 drivers
v0x5c7c32ef9a60_0 .net "in_b", 0 0, L_0x5c7c33111c30;  alias, 1 drivers
v0x5c7c32ef9b50_0 .net "out", 0 0, L_0x5c7c33111ce0;  alias, 1 drivers
S_0x5c7c32efa100 .scope module, "xor_gate" "Xor" 4 8, 8 2 0, S_0x5c7c32ef8b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f03ef0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32f03f90_0 .net "in_b", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32f04050_0 .net "out", 0 0, L_0x5c7c33112950;  alias, 1 drivers
v0x5c7c32f040f0_0 .net "temp_a_and_out", 0 0, L_0x5c7c33111ef0;  1 drivers
v0x5c7c32f042a0_0 .net "temp_a_out", 0 0, L_0x5c7c33111d90;  1 drivers
v0x5c7c32f04340_0 .net "temp_b_and_out", 0 0, L_0x5c7c33112100;  1 drivers
v0x5c7c32f044f0_0 .net "temp_b_out", 0 0, L_0x5c7c33111fa0;  1 drivers
S_0x5c7c32efa2e0 .scope module, "and_gate" "And" 8 10, 5 2 0, S_0x5c7c32efa100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32efb3d0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32efb470_0 .net "in_b", 0 0, L_0x5c7c33111d90;  alias, 1 drivers
v0x5c7c32efb560_0 .net "out", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
v0x5c7c32efb680_0 .net "temp_out", 0 0, L_0x5c7c33111e40;  1 drivers
S_0x5c7c32efa550 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32efa2e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33111e40 .functor NAND 1, L_0x5c7c33112b10, L_0x5c7c33111d90, C4<1>, C4<1>;
v0x5c7c32efa7c0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32efa8d0_0 .net "in_b", 0 0, L_0x5c7c33111d90;  alias, 1 drivers
v0x5c7c32efa990_0 .net "out", 0 0, L_0x5c7c33111e40;  alias, 1 drivers
S_0x5c7c32efaab0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32efa2e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32efb220_0 .net "in_a", 0 0, L_0x5c7c33111e40;  alias, 1 drivers
v0x5c7c32efb2c0_0 .net "out", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
S_0x5c7c32efacd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32efaab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33111ef0 .functor NAND 1, L_0x5c7c33111e40, L_0x5c7c33111e40, C4<1>, C4<1>;
v0x5c7c32efaf40_0 .net "in_a", 0 0, L_0x5c7c33111e40;  alias, 1 drivers
v0x5c7c32efb030_0 .net "in_b", 0 0, L_0x5c7c33111e40;  alias, 1 drivers
v0x5c7c32efb120_0 .net "out", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
S_0x5c7c32efb740 .scope module, "and_gate2" "And" 8 14, 5 2 0, S_0x5c7c32efa100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32efc770_0 .net "in_a", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32efc810_0 .net "in_b", 0 0, L_0x5c7c33111fa0;  alias, 1 drivers
v0x5c7c32efc900_0 .net "out", 0 0, L_0x5c7c33112100;  alias, 1 drivers
v0x5c7c32efca20_0 .net "temp_out", 0 0, L_0x5c7c33112050;  1 drivers
S_0x5c7c32efb920 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32efb740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112050 .functor NAND 1, L_0x5c7c33112be0, L_0x5c7c33111fa0, C4<1>, C4<1>;
v0x5c7c32efbb90_0 .net "in_a", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32efbca0_0 .net "in_b", 0 0, L_0x5c7c33111fa0;  alias, 1 drivers
v0x5c7c32efbd60_0 .net "out", 0 0, L_0x5c7c33112050;  alias, 1 drivers
S_0x5c7c32efbe80 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32efb740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32efc5c0_0 .net "in_a", 0 0, L_0x5c7c33112050;  alias, 1 drivers
v0x5c7c32efc660_0 .net "out", 0 0, L_0x5c7c33112100;  alias, 1 drivers
S_0x5c7c32efc0a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32efbe80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112100 .functor NAND 1, L_0x5c7c33112050, L_0x5c7c33112050, C4<1>, C4<1>;
v0x5c7c32efc310_0 .net "in_a", 0 0, L_0x5c7c33112050;  alias, 1 drivers
v0x5c7c32efc3d0_0 .net "in_b", 0 0, L_0x5c7c33112050;  alias, 1 drivers
v0x5c7c32efc4c0_0 .net "out", 0 0, L_0x5c7c33112100;  alias, 1 drivers
S_0x5c7c32efcb70 .scope module, "not_gate" "Not" 8 9, 7 3 0, S_0x5c7c32efa100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32efd2b0_0 .net "in_a", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32efd350_0 .net "out", 0 0, L_0x5c7c33111d90;  alias, 1 drivers
S_0x5c7c32efcd40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32efcb70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33111d90 .functor NAND 1, L_0x5c7c33112be0, L_0x5c7c33112be0, C4<1>, C4<1>;
v0x5c7c32efcf90_0 .net "in_a", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32efd0e0_0 .net "in_b", 0 0, L_0x5c7c33112be0;  alias, 1 drivers
v0x5c7c32efd1a0_0 .net "out", 0 0, L_0x5c7c33111d90;  alias, 1 drivers
S_0x5c7c32efd450 .scope module, "not_gate2" "Not" 8 13, 7 3 0, S_0x5c7c32efa100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32efdbd0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32efdc70_0 .net "out", 0 0, L_0x5c7c33111fa0;  alias, 1 drivers
S_0x5c7c32efd670 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32efd450;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33111fa0 .functor NAND 1, L_0x5c7c33112b10, L_0x5c7c33112b10, C4<1>, C4<1>;
v0x5c7c32efd8e0_0 .net "in_a", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32efda30_0 .net "in_b", 0 0, L_0x5c7c33112b10;  alias, 1 drivers
v0x5c7c32efdaf0_0 .net "out", 0 0, L_0x5c7c33111fa0;  alias, 1 drivers
S_0x5c7c32efdd70 .scope module, "or_gate" "Or" 8 17, 9 3 0, S_0x5c7c32efa100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f03840_0 .net "branch1_out", 0 0, L_0x5c7c33112310;  1 drivers
v0x5c7c32f03970_0 .net "branch2_out", 0 0, L_0x5c7c33112630;  1 drivers
v0x5c7c32f03ac0_0 .net "in_a", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
v0x5c7c32f03b90_0 .net "in_b", 0 0, L_0x5c7c33112100;  alias, 1 drivers
v0x5c7c32f03c30_0 .net "out", 0 0, L_0x5c7c33112950;  alias, 1 drivers
v0x5c7c32f03cd0_0 .net "temp1_out", 0 0, L_0x5c7c33112260;  1 drivers
v0x5c7c32f03d70_0 .net "temp2_out", 0 0, L_0x5c7c33112580;  1 drivers
v0x5c7c32f03e10_0 .net "temp3_out", 0 0, L_0x5c7c331128a0;  1 drivers
S_0x5c7c32efdff0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32efdd70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32eff080_0 .net "in_a", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
v0x5c7c32eff120_0 .net "in_b", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
v0x5c7c32eff1e0_0 .net "out", 0 0, L_0x5c7c33112260;  alias, 1 drivers
v0x5c7c32eff300_0 .net "temp_out", 0 0, L_0x5c7c331121b0;  1 drivers
S_0x5c7c32efe260 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32efdff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331121b0 .functor NAND 1, L_0x5c7c33111ef0, L_0x5c7c33111ef0, C4<1>, C4<1>;
v0x5c7c32efe4d0_0 .net "in_a", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
v0x5c7c32efe590_0 .net "in_b", 0 0, L_0x5c7c33111ef0;  alias, 1 drivers
v0x5c7c32efe6e0_0 .net "out", 0 0, L_0x5c7c331121b0;  alias, 1 drivers
S_0x5c7c32efe7e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32efdff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32efeed0_0 .net "in_a", 0 0, L_0x5c7c331121b0;  alias, 1 drivers
v0x5c7c32efef70_0 .net "out", 0 0, L_0x5c7c33112260;  alias, 1 drivers
S_0x5c7c32efe9b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32efe7e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112260 .functor NAND 1, L_0x5c7c331121b0, L_0x5c7c331121b0, C4<1>, C4<1>;
v0x5c7c32efec20_0 .net "in_a", 0 0, L_0x5c7c331121b0;  alias, 1 drivers
v0x5c7c32efece0_0 .net "in_b", 0 0, L_0x5c7c331121b0;  alias, 1 drivers
v0x5c7c32efedd0_0 .net "out", 0 0, L_0x5c7c33112260;  alias, 1 drivers
S_0x5c7c32eff470 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32efdd70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f004a0_0 .net "in_a", 0 0, L_0x5c7c33112100;  alias, 1 drivers
v0x5c7c32f00540_0 .net "in_b", 0 0, L_0x5c7c33112100;  alias, 1 drivers
v0x5c7c32f00600_0 .net "out", 0 0, L_0x5c7c33112580;  alias, 1 drivers
v0x5c7c32f00720_0 .net "temp_out", 0 0, L_0x5c7c331124d0;  1 drivers
S_0x5c7c32eff650 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32eff470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331124d0 .functor NAND 1, L_0x5c7c33112100, L_0x5c7c33112100, C4<1>, C4<1>;
v0x5c7c32eff8c0_0 .net "in_a", 0 0, L_0x5c7c33112100;  alias, 1 drivers
v0x5c7c32eff980_0 .net "in_b", 0 0, L_0x5c7c33112100;  alias, 1 drivers
v0x5c7c32effad0_0 .net "out", 0 0, L_0x5c7c331124d0;  alias, 1 drivers
S_0x5c7c32effbd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32eff470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f002f0_0 .net "in_a", 0 0, L_0x5c7c331124d0;  alias, 1 drivers
v0x5c7c32f00390_0 .net "out", 0 0, L_0x5c7c33112580;  alias, 1 drivers
S_0x5c7c32effda0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32effbd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112580 .functor NAND 1, L_0x5c7c331124d0, L_0x5c7c331124d0, C4<1>, C4<1>;
v0x5c7c32f00010_0 .net "in_a", 0 0, L_0x5c7c331124d0;  alias, 1 drivers
v0x5c7c32f00100_0 .net "in_b", 0 0, L_0x5c7c331124d0;  alias, 1 drivers
v0x5c7c32f001f0_0 .net "out", 0 0, L_0x5c7c33112580;  alias, 1 drivers
S_0x5c7c32f00890 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32efdd70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f018d0_0 .net "in_a", 0 0, L_0x5c7c33112310;  alias, 1 drivers
v0x5c7c32f019a0_0 .net "in_b", 0 0, L_0x5c7c33112630;  alias, 1 drivers
v0x5c7c32f01a70_0 .net "out", 0 0, L_0x5c7c331128a0;  alias, 1 drivers
v0x5c7c32f01b90_0 .net "temp_out", 0 0, L_0x5c7c331127f0;  1 drivers
S_0x5c7c32f00a70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f00890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331127f0 .functor NAND 1, L_0x5c7c33112310, L_0x5c7c33112630, C4<1>, C4<1>;
v0x5c7c32f00cc0_0 .net "in_a", 0 0, L_0x5c7c33112310;  alias, 1 drivers
v0x5c7c32f00da0_0 .net "in_b", 0 0, L_0x5c7c33112630;  alias, 1 drivers
v0x5c7c32f00e60_0 .net "out", 0 0, L_0x5c7c331127f0;  alias, 1 drivers
S_0x5c7c32f00fb0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f00890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f01720_0 .net "in_a", 0 0, L_0x5c7c331127f0;  alias, 1 drivers
v0x5c7c32f017c0_0 .net "out", 0 0, L_0x5c7c331128a0;  alias, 1 drivers
S_0x5c7c32f011d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f00fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331128a0 .functor NAND 1, L_0x5c7c331127f0, L_0x5c7c331127f0, C4<1>, C4<1>;
v0x5c7c32f01440_0 .net "in_a", 0 0, L_0x5c7c331127f0;  alias, 1 drivers
v0x5c7c32f01530_0 .net "in_b", 0 0, L_0x5c7c331127f0;  alias, 1 drivers
v0x5c7c32f01620_0 .net "out", 0 0, L_0x5c7c331128a0;  alias, 1 drivers
S_0x5c7c32f01ce0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32efdd70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f02410_0 .net "in_a", 0 0, L_0x5c7c33112260;  alias, 1 drivers
v0x5c7c32f024b0_0 .net "out", 0 0, L_0x5c7c33112310;  alias, 1 drivers
S_0x5c7c32f01eb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f01ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112310 .functor NAND 1, L_0x5c7c33112260, L_0x5c7c33112260, C4<1>, C4<1>;
v0x5c7c32f02120_0 .net "in_a", 0 0, L_0x5c7c33112260;  alias, 1 drivers
v0x5c7c32f021e0_0 .net "in_b", 0 0, L_0x5c7c33112260;  alias, 1 drivers
v0x5c7c32f02330_0 .net "out", 0 0, L_0x5c7c33112310;  alias, 1 drivers
S_0x5c7c32f025b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32efdd70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f02d80_0 .net "in_a", 0 0, L_0x5c7c33112580;  alias, 1 drivers
v0x5c7c32f02e20_0 .net "out", 0 0, L_0x5c7c33112630;  alias, 1 drivers
S_0x5c7c32f02820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f025b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112630 .functor NAND 1, L_0x5c7c33112580, L_0x5c7c33112580, C4<1>, C4<1>;
v0x5c7c32f02a90_0 .net "in_a", 0 0, L_0x5c7c33112580;  alias, 1 drivers
v0x5c7c32f02b50_0 .net "in_b", 0 0, L_0x5c7c33112580;  alias, 1 drivers
v0x5c7c32f02ca0_0 .net "out", 0 0, L_0x5c7c33112630;  alias, 1 drivers
S_0x5c7c32f02f20 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32efdd70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f036c0_0 .net "in_a", 0 0, L_0x5c7c331128a0;  alias, 1 drivers
v0x5c7c32f03760_0 .net "out", 0 0, L_0x5c7c33112950;  alias, 1 drivers
S_0x5c7c32f03140 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f02f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33112950 .functor NAND 1, L_0x5c7c331128a0, L_0x5c7c331128a0, C4<1>, C4<1>;
v0x5c7c32f033b0_0 .net "in_a", 0 0, L_0x5c7c331128a0;  alias, 1 drivers
v0x5c7c32f03470_0 .net "in_b", 0 0, L_0x5c7c331128a0;  alias, 1 drivers
v0x5c7c32f035c0_0 .net "out", 0 0, L_0x5c7c33112950;  alias, 1 drivers
S_0x5c7c32d01140 .scope module, "And16" "And16" 10 2;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "in_a";
    .port_info 1 /INPUT 16 "in_b";
    .port_info 2 /OUTPUT 16 "out";
o0x7d2eeb8620a8 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c32f10190_0 .net "in_a", 15 0, o0x7d2eeb8620a8;  0 drivers
o0x7d2eeb8620d8 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c32f10270_0 .net "in_b", 15 0, o0x7d2eeb8620d8;  0 drivers
v0x5c7c32f10350_0 .net "out", 15 0, L_0x5c7c3313d1d0;  1 drivers
v0x5c7c32f10450_0 .net/s "temp_out", 15 0, L_0x5c7c33139d50;  1 drivers
L_0x5c7c33136af0 .part o0x7d2eeb8620a8, 0, 1;
L_0x5c7c33136b90 .part o0x7d2eeb8620d8, 0, 1;
L_0x5c7c33136d30 .part o0x7d2eeb8620a8, 1, 1;
L_0x5c7c33136e20 .part o0x7d2eeb8620d8, 1, 1;
L_0x5c7c33137000 .part o0x7d2eeb8620a8, 2, 1;
L_0x5c7c331370f0 .part o0x7d2eeb8620d8, 2, 1;
L_0x5c7c33137290 .part o0x7d2eeb8620a8, 3, 1;
L_0x5c7c33137380 .part o0x7d2eeb8620d8, 3, 1;
L_0x5c7c331374e0 .part o0x7d2eeb8620a8, 4, 1;
L_0x5c7c33137580 .part o0x7d2eeb8620d8, 4, 1;
L_0x5c7c33137770 .part o0x7d2eeb8620a8, 5, 1;
L_0x5c7c33137810 .part o0x7d2eeb8620d8, 5, 1;
L_0x5c7c33137a10 .part o0x7d2eeb8620a8, 6, 1;
L_0x5c7c33137b00 .part o0x7d2eeb8620d8, 6, 1;
L_0x5c7c33137ca0 .part o0x7d2eeb8620a8, 7, 1;
L_0x5c7c33137d90 .part o0x7d2eeb8620d8, 7, 1;
L_0x5c7c33137fb0 .part o0x7d2eeb8620a8, 8, 1;
L_0x5c7c331380a0 .part o0x7d2eeb8620d8, 8, 1;
L_0x5c7c331382d0 .part o0x7d2eeb8620a8, 9, 1;
L_0x5c7c331383c0 .part o0x7d2eeb8620d8, 9, 1;
L_0x5c7c33138190 .part o0x7d2eeb8620a8, 10, 1;
L_0x5c7c33138650 .part o0x7d2eeb8620d8, 10, 1;
L_0x5c7c331388a0 .part o0x7d2eeb8620a8, 11, 1;
L_0x5c7c33138990 .part o0x7d2eeb8620d8, 11, 1;
L_0x5c7c33138bf0 .part o0x7d2eeb8620a8, 12, 1;
L_0x5c7c33138ce0 .part o0x7d2eeb8620d8, 12, 1;
L_0x5c7c33138f50 .part o0x7d2eeb8620a8, 13, 1;
L_0x5c7c33139040 .part o0x7d2eeb8620d8, 13, 1;
L_0x5c7c331392c0 .part o0x7d2eeb8620a8, 14, 1;
L_0x5c7c331393b0 .part o0x7d2eeb8620d8, 14, 1;
L_0x5c7c33139640 .part o0x7d2eeb8620a8, 15, 1;
L_0x5c7c33139940 .part o0x7d2eeb8620d8, 15, 1;
LS_0x5c7c33139d50_0_0 .concat8 [ 1 1 1 1], L_0x5c7c32de2bf0, L_0x5c7c33136c30, L_0x5c7c33136f90, L_0x5c7c33137220;
LS_0x5c7c33139d50_0_4 .concat8 [ 1 1 1 1], L_0x5c7c33137470, L_0x5c7c331376d0, L_0x5c7c33137970, L_0x5c7c33137900;
LS_0x5c7c33139d50_0_8 .concat8 [ 1 1 1 1], L_0x5c7c33137f10, L_0x5c7c33138230, L_0x5c7c33138560, L_0x5c7c33138800;
LS_0x5c7c33139d50_0_12 .concat8 [ 1 1 1 1], L_0x5c7c33138b50, L_0x5c7c33138eb0, L_0x5c7c33139220, L_0x5c7c331395a0;
L_0x5c7c33139d50 .concat8 [ 4 4 4 4], LS_0x5c7c33139d50_0_0, LS_0x5c7c33139d50_0_4, LS_0x5c7c33139d50_0_8, LS_0x5c7c33139d50_0_12;
S_0x5c7c32f05990 .scope module, "nand_gate0" "Nand" 10 5, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32de2bf0 .functor NAND 1, L_0x5c7c33136af0, L_0x5c7c33136b90, C4<1>, C4<1>;
v0x5c7c32f05b40_0 .net "in_a", 0 0, L_0x5c7c33136af0;  1 drivers
v0x5c7c32f05c20_0 .net "in_b", 0 0, L_0x5c7c33136b90;  1 drivers
v0x5c7c32f05ce0_0 .net "out", 0 0, L_0x5c7c32de2bf0;  1 drivers
S_0x5c7c32f05e00 .scope module, "nand_gate1" "Nand" 10 6, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33136c30 .functor NAND 1, L_0x5c7c33136d30, L_0x5c7c33136e20, C4<1>, C4<1>;
v0x5c7c32f05f90_0 .net "in_a", 0 0, L_0x5c7c33136d30;  1 drivers
v0x5c7c32f06070_0 .net "in_b", 0 0, L_0x5c7c33136e20;  1 drivers
v0x5c7c32f06130_0 .net "out", 0 0, L_0x5c7c33136c30;  1 drivers
S_0x5c7c32f06280 .scope module, "nand_gate10" "Nand" 10 15, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33138560 .functor NAND 1, L_0x5c7c33138190, L_0x5c7c33138650, C4<1>, C4<1>;
v0x5c7c32f064e0_0 .net "in_a", 0 0, L_0x5c7c33138190;  1 drivers
v0x5c7c32f065a0_0 .net "in_b", 0 0, L_0x5c7c33138650;  1 drivers
v0x5c7c32f06660_0 .net "out", 0 0, L_0x5c7c33138560;  1 drivers
S_0x5c7c32f067b0 .scope module, "nand_gate11" "Nand" 10 16, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33138800 .functor NAND 1, L_0x5c7c331388a0, L_0x5c7c33138990, C4<1>, C4<1>;
v0x5c7c32f069e0_0 .net "in_a", 0 0, L_0x5c7c331388a0;  1 drivers
v0x5c7c32f06ac0_0 .net "in_b", 0 0, L_0x5c7c33138990;  1 drivers
v0x5c7c32f06b80_0 .net "out", 0 0, L_0x5c7c33138800;  1 drivers
S_0x5c7c32f06cd0 .scope module, "nand_gate12" "Nand" 10 17, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33138b50 .functor NAND 1, L_0x5c7c33138bf0, L_0x5c7c33138ce0, C4<1>, C4<1>;
v0x5c7c32f06f50_0 .net "in_a", 0 0, L_0x5c7c33138bf0;  1 drivers
v0x5c7c32f07030_0 .net "in_b", 0 0, L_0x5c7c33138ce0;  1 drivers
v0x5c7c32f070f0_0 .net "out", 0 0, L_0x5c7c33138b50;  1 drivers
S_0x5c7c32f07210 .scope module, "nand_gate13" "Nand" 10 18, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33138eb0 .functor NAND 1, L_0x5c7c33138f50, L_0x5c7c33139040, C4<1>, C4<1>;
v0x5c7c32f07440_0 .net "in_a", 0 0, L_0x5c7c33138f50;  1 drivers
v0x5c7c32f07520_0 .net "in_b", 0 0, L_0x5c7c33139040;  1 drivers
v0x5c7c32f075e0_0 .net "out", 0 0, L_0x5c7c33138eb0;  1 drivers
S_0x5c7c32f07730 .scope module, "nand_gate14" "Nand" 10 19, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33139220 .functor NAND 1, L_0x5c7c331392c0, L_0x5c7c331393b0, C4<1>, C4<1>;
v0x5c7c32f07960_0 .net "in_a", 0 0, L_0x5c7c331392c0;  1 drivers
v0x5c7c32f07a40_0 .net "in_b", 0 0, L_0x5c7c331393b0;  1 drivers
v0x5c7c32f07b00_0 .net "out", 0 0, L_0x5c7c33139220;  1 drivers
S_0x5c7c32f07c50 .scope module, "nand_gate15" "Nand" 10 20, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331395a0 .functor NAND 1, L_0x5c7c33139640, L_0x5c7c33139940, C4<1>, C4<1>;
v0x5c7c32f07e80_0 .net "in_a", 0 0, L_0x5c7c33139640;  1 drivers
v0x5c7c32f07f60_0 .net "in_b", 0 0, L_0x5c7c33139940;  1 drivers
v0x5c7c32f08020_0 .net "out", 0 0, L_0x5c7c331395a0;  1 drivers
S_0x5c7c32f08170 .scope module, "nand_gate2" "Nand" 10 7, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33136f90 .functor NAND 1, L_0x5c7c33137000, L_0x5c7c331370f0, C4<1>, C4<1>;
v0x5c7c32f08350_0 .net "in_a", 0 0, L_0x5c7c33137000;  1 drivers
v0x5c7c32f08430_0 .net "in_b", 0 0, L_0x5c7c331370f0;  1 drivers
v0x5c7c32f084f0_0 .net "out", 0 0, L_0x5c7c33136f90;  1 drivers
S_0x5c7c32f08640 .scope module, "nand_gate3" "Nand" 10 8, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33137220 .functor NAND 1, L_0x5c7c33137290, L_0x5c7c33137380, C4<1>, C4<1>;
v0x5c7c32f08870_0 .net "in_a", 0 0, L_0x5c7c33137290;  1 drivers
v0x5c7c32f08950_0 .net "in_b", 0 0, L_0x5c7c33137380;  1 drivers
v0x5c7c32f08a10_0 .net "out", 0 0, L_0x5c7c33137220;  1 drivers
S_0x5c7c32f08b60 .scope module, "nand_gate4" "Nand" 10 9, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33137470 .functor NAND 1, L_0x5c7c331374e0, L_0x5c7c33137580, C4<1>, C4<1>;
v0x5c7c32f08d90_0 .net "in_a", 0 0, L_0x5c7c331374e0;  1 drivers
v0x5c7c32f08e70_0 .net "in_b", 0 0, L_0x5c7c33137580;  1 drivers
v0x5c7c32f08f30_0 .net "out", 0 0, L_0x5c7c33137470;  1 drivers
S_0x5c7c32f09080 .scope module, "nand_gate5" "Nand" 10 10, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331376d0 .functor NAND 1, L_0x5c7c33137770, L_0x5c7c33137810, C4<1>, C4<1>;
v0x5c7c32f092b0_0 .net "in_a", 0 0, L_0x5c7c33137770;  1 drivers
v0x5c7c32f09390_0 .net "in_b", 0 0, L_0x5c7c33137810;  1 drivers
v0x5c7c32f09450_0 .net "out", 0 0, L_0x5c7c331376d0;  1 drivers
S_0x5c7c32f095a0 .scope module, "nand_gate6" "Nand" 10 11, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33137970 .functor NAND 1, L_0x5c7c33137a10, L_0x5c7c33137b00, C4<1>, C4<1>;
v0x5c7c32f097d0_0 .net "in_a", 0 0, L_0x5c7c33137a10;  1 drivers
v0x5c7c32f098b0_0 .net "in_b", 0 0, L_0x5c7c33137b00;  1 drivers
v0x5c7c32f09970_0 .net "out", 0 0, L_0x5c7c33137970;  1 drivers
S_0x5c7c32f09ac0 .scope module, "nand_gate7" "Nand" 10 12, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33137900 .functor NAND 1, L_0x5c7c33137ca0, L_0x5c7c33137d90, C4<1>, C4<1>;
v0x5c7c32f09cf0_0 .net "in_a", 0 0, L_0x5c7c33137ca0;  1 drivers
v0x5c7c32f09dd0_0 .net "in_b", 0 0, L_0x5c7c33137d90;  1 drivers
v0x5c7c32f09e90_0 .net "out", 0 0, L_0x5c7c33137900;  1 drivers
S_0x5c7c32f09fe0 .scope module, "nand_gate8" "Nand" 10 13, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33137f10 .functor NAND 1, L_0x5c7c33137fb0, L_0x5c7c331380a0, C4<1>, C4<1>;
v0x5c7c32f0a210_0 .net "in_a", 0 0, L_0x5c7c33137fb0;  1 drivers
v0x5c7c32f0a2f0_0 .net "in_b", 0 0, L_0x5c7c331380a0;  1 drivers
v0x5c7c32f0a3b0_0 .net "out", 0 0, L_0x5c7c33137f10;  1 drivers
S_0x5c7c32f0a500 .scope module, "nand_gate9" "Nand" 10 14, 6 1 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33138230 .functor NAND 1, L_0x5c7c331382d0, L_0x5c7c331383c0, C4<1>, C4<1>;
v0x5c7c32f0a730_0 .net "in_a", 0 0, L_0x5c7c331382d0;  1 drivers
v0x5c7c32f0a810_0 .net "in_b", 0 0, L_0x5c7c331383c0;  1 drivers
v0x5c7c32f0a8d0_0 .net "out", 0 0, L_0x5c7c33138230;  1 drivers
S_0x5c7c32f0aa20 .scope module, "not16_gate" "Not16" 10 22, 11 3 0, S_0x5c7c32d01140;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "in_a";
    .port_info 1 /OUTPUT 16 "out";
v0x5c7c32f0ff70_0 .net "in_a", 15 0, L_0x5c7c33139d50;  alias, 1 drivers
v0x5c7c32f10050_0 .net "out", 15 0, L_0x5c7c3313d1d0;  alias, 1 drivers
L_0x5c7c3313a3b0 .part L_0x5c7c33139d50, 0, 1;
L_0x5c7c3313a4a0 .part L_0x5c7c33139d50, 0, 1;
L_0x5c7c3313a600 .part L_0x5c7c33139d50, 1, 1;
L_0x5c7c3313a6a0 .part L_0x5c7c33139d50, 1, 1;
L_0x5c7c3313a800 .part L_0x5c7c33139d50, 2, 1;
L_0x5c7c3313a8f0 .part L_0x5c7c33139d50, 2, 1;
L_0x5c7c3313aa90 .part L_0x5c7c33139d50, 3, 1;
L_0x5c7c3313ab80 .part L_0x5c7c33139d50, 3, 1;
L_0x5c7c3313ad30 .part L_0x5c7c33139d50, 4, 1;
L_0x5c7c3313ae20 .part L_0x5c7c33139d50, 4, 1;
L_0x5c7c3313afe0 .part L_0x5c7c33139d50, 5, 1;
L_0x5c7c3313b080 .part L_0x5c7c33139d50, 5, 1;
L_0x5c7c3313b250 .part L_0x5c7c33139d50, 6, 1;
L_0x5c7c3313b340 .part L_0x5c7c33139d50, 6, 1;
L_0x5c7c3313b6c0 .part L_0x5c7c33139d50, 7, 1;
L_0x5c7c3313b7b0 .part L_0x5c7c33139d50, 7, 1;
L_0x5c7c3313b9a0 .part L_0x5c7c33139d50, 8, 1;
L_0x5c7c3313ba90 .part L_0x5c7c33139d50, 8, 1;
L_0x5c7c3313bc90 .part L_0x5c7c33139d50, 9, 1;
L_0x5c7c3313bd80 .part L_0x5c7c33139d50, 9, 1;
L_0x5c7c3313bb80 .part L_0x5c7c33139d50, 10, 1;
L_0x5c7c3313bfe0 .part L_0x5c7c33139d50, 10, 1;
L_0x5c7c3313c200 .part L_0x5c7c33139d50, 11, 1;
L_0x5c7c3313c2f0 .part L_0x5c7c33139d50, 11, 1;
L_0x5c7c3313c520 .part L_0x5c7c33139d50, 12, 1;
L_0x5c7c3313c610 .part L_0x5c7c33139d50, 12, 1;
L_0x5c7c3313c850 .part L_0x5c7c33139d50, 13, 1;
L_0x5c7c3313c940 .part L_0x5c7c33139d50, 13, 1;
L_0x5c7c3313cb90 .part L_0x5c7c33139d50, 14, 1;
L_0x5c7c3313cc80 .part L_0x5c7c33139d50, 14, 1;
L_0x5c7c3313cee0 .part L_0x5c7c33139d50, 15, 1;
L_0x5c7c3313cfd0 .part L_0x5c7c33139d50, 15, 1;
LS_0x5c7c3313d1d0_0_0 .concat8 [ 1 1 1 1], L_0x5c7c3313a340, L_0x5c7c3313a590, L_0x5c7c3313a790, L_0x5c7c3313aa20;
LS_0x5c7c3313d1d0_0_4 .concat8 [ 1 1 1 1], L_0x5c7c3313acc0, L_0x5c7c3313af70, L_0x5c7c3313b1e0, L_0x5c7c3313b170;
LS_0x5c7c3313d1d0_0_8 .concat8 [ 1 1 1 1], L_0x5c7c3313b930, L_0x5c7c3313bc20, L_0x5c7c3313bf20, L_0x5c7c3313c190;
LS_0x5c7c3313d1d0_0_12 .concat8 [ 1 1 1 1], L_0x5c7c3313c4b0, L_0x5c7c3313c7e0, L_0x5c7c3313cb20, L_0x5c7c3313ce70;
L_0x5c7c3313d1d0 .concat8 [ 4 4 4 4], LS_0x5c7c3313d1d0_0_0, LS_0x5c7c3313d1d0_0_4, LS_0x5c7c3313d1d0_0_8, LS_0x5c7c3313d1d0_0_12;
S_0x5c7c32f0ad50 .scope module, "nand_gate0" "Nand" 11 4, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313a340 .functor NAND 1, L_0x5c7c3313a3b0, L_0x5c7c3313a4a0, C4<1>, C4<1>;
v0x5c7c32f0afc0_0 .net "in_a", 0 0, L_0x5c7c3313a3b0;  1 drivers
v0x5c7c32f0b0a0_0 .net "in_b", 0 0, L_0x5c7c3313a4a0;  1 drivers
v0x5c7c32f0b160_0 .net "out", 0 0, L_0x5c7c3313a340;  1 drivers
S_0x5c7c32f0b2b0 .scope module, "nand_gate1" "Nand" 11 5, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313a590 .functor NAND 1, L_0x5c7c3313a600, L_0x5c7c3313a6a0, C4<1>, C4<1>;
v0x5c7c32f0b4e0_0 .net "in_a", 0 0, L_0x5c7c3313a600;  1 drivers
v0x5c7c32f0b5c0_0 .net "in_b", 0 0, L_0x5c7c3313a6a0;  1 drivers
v0x5c7c32f0b680_0 .net "out", 0 0, L_0x5c7c3313a590;  1 drivers
S_0x5c7c32f0b7d0 .scope module, "nand_gate10" "Nand" 11 14, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313bf20 .functor NAND 1, L_0x5c7c3313bb80, L_0x5c7c3313bfe0, C4<1>, C4<1>;
v0x5c7c32f0ba30_0 .net "in_a", 0 0, L_0x5c7c3313bb80;  1 drivers
v0x5c7c32f0baf0_0 .net "in_b", 0 0, L_0x5c7c3313bfe0;  1 drivers
v0x5c7c32f0bbb0_0 .net "out", 0 0, L_0x5c7c3313bf20;  1 drivers
S_0x5c7c32f0bd00 .scope module, "nand_gate11" "Nand" 11 15, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313c190 .functor NAND 1, L_0x5c7c3313c200, L_0x5c7c3313c2f0, C4<1>, C4<1>;
v0x5c7c32f0bf30_0 .net "in_a", 0 0, L_0x5c7c3313c200;  1 drivers
v0x5c7c32f0c010_0 .net "in_b", 0 0, L_0x5c7c3313c2f0;  1 drivers
v0x5c7c32f0c0d0_0 .net "out", 0 0, L_0x5c7c3313c190;  1 drivers
S_0x5c7c32f0c220 .scope module, "nand_gate12" "Nand" 11 16, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313c4b0 .functor NAND 1, L_0x5c7c3313c520, L_0x5c7c3313c610, C4<1>, C4<1>;
v0x5c7c32f0c4a0_0 .net "in_a", 0 0, L_0x5c7c3313c520;  1 drivers
v0x5c7c32f0c580_0 .net "in_b", 0 0, L_0x5c7c3313c610;  1 drivers
v0x5c7c32f0c640_0 .net "out", 0 0, L_0x5c7c3313c4b0;  1 drivers
S_0x5c7c32f0c760 .scope module, "nand_gate13" "Nand" 11 17, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313c7e0 .functor NAND 1, L_0x5c7c3313c850, L_0x5c7c3313c940, C4<1>, C4<1>;
v0x5c7c32f0c990_0 .net "in_a", 0 0, L_0x5c7c3313c850;  1 drivers
v0x5c7c32f0ca70_0 .net "in_b", 0 0, L_0x5c7c3313c940;  1 drivers
v0x5c7c32f0cb30_0 .net "out", 0 0, L_0x5c7c3313c7e0;  1 drivers
S_0x5c7c32f0cc80 .scope module, "nand_gate14" "Nand" 11 18, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313cb20 .functor NAND 1, L_0x5c7c3313cb90, L_0x5c7c3313cc80, C4<1>, C4<1>;
v0x5c7c32f0ceb0_0 .net "in_a", 0 0, L_0x5c7c3313cb90;  1 drivers
v0x5c7c32f0cf90_0 .net "in_b", 0 0, L_0x5c7c3313cc80;  1 drivers
v0x5c7c32f0d050_0 .net "out", 0 0, L_0x5c7c3313cb20;  1 drivers
S_0x5c7c32f0d1a0 .scope module, "nand_gate15" "Nand" 11 19, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313ce70 .functor NAND 1, L_0x5c7c3313cee0, L_0x5c7c3313cfd0, C4<1>, C4<1>;
v0x5c7c32f0d3d0_0 .net "in_a", 0 0, L_0x5c7c3313cee0;  1 drivers
v0x5c7c32f0d4b0_0 .net "in_b", 0 0, L_0x5c7c3313cfd0;  1 drivers
v0x5c7c32f0d570_0 .net "out", 0 0, L_0x5c7c3313ce70;  1 drivers
S_0x5c7c32f0d6c0 .scope module, "nand_gate2" "Nand" 11 6, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313a790 .functor NAND 1, L_0x5c7c3313a800, L_0x5c7c3313a8f0, C4<1>, C4<1>;
v0x5c7c32f0d8a0_0 .net "in_a", 0 0, L_0x5c7c3313a800;  1 drivers
v0x5c7c32f0d980_0 .net "in_b", 0 0, L_0x5c7c3313a8f0;  1 drivers
v0x5c7c32f0da40_0 .net "out", 0 0, L_0x5c7c3313a790;  1 drivers
S_0x5c7c32f0db90 .scope module, "nand_gate3" "Nand" 11 7, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313aa20 .functor NAND 1, L_0x5c7c3313aa90, L_0x5c7c3313ab80, C4<1>, C4<1>;
v0x5c7c32f0ddc0_0 .net "in_a", 0 0, L_0x5c7c3313aa90;  1 drivers
v0x5c7c32f0dea0_0 .net "in_b", 0 0, L_0x5c7c3313ab80;  1 drivers
v0x5c7c32f0df60_0 .net "out", 0 0, L_0x5c7c3313aa20;  1 drivers
S_0x5c7c32f0e0b0 .scope module, "nand_gate4" "Nand" 11 8, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313acc0 .functor NAND 1, L_0x5c7c3313ad30, L_0x5c7c3313ae20, C4<1>, C4<1>;
v0x5c7c32f0e2e0_0 .net "in_a", 0 0, L_0x5c7c3313ad30;  1 drivers
v0x5c7c32f0e3c0_0 .net "in_b", 0 0, L_0x5c7c3313ae20;  1 drivers
v0x5c7c32f0e480_0 .net "out", 0 0, L_0x5c7c3313acc0;  1 drivers
S_0x5c7c32f0e5d0 .scope module, "nand_gate5" "Nand" 11 9, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313af70 .functor NAND 1, L_0x5c7c3313afe0, L_0x5c7c3313b080, C4<1>, C4<1>;
v0x5c7c32f0e800_0 .net "in_a", 0 0, L_0x5c7c3313afe0;  1 drivers
v0x5c7c32f0e8e0_0 .net "in_b", 0 0, L_0x5c7c3313b080;  1 drivers
v0x5c7c32f0e9a0_0 .net "out", 0 0, L_0x5c7c3313af70;  1 drivers
S_0x5c7c32f0eaf0 .scope module, "nand_gate6" "Nand" 11 10, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313b1e0 .functor NAND 1, L_0x5c7c3313b250, L_0x5c7c3313b340, C4<1>, C4<1>;
v0x5c7c32f0ed20_0 .net "in_a", 0 0, L_0x5c7c3313b250;  1 drivers
v0x5c7c32f0ee00_0 .net "in_b", 0 0, L_0x5c7c3313b340;  1 drivers
v0x5c7c32f0eec0_0 .net "out", 0 0, L_0x5c7c3313b1e0;  1 drivers
S_0x5c7c32f0f010 .scope module, "nand_gate7" "Nand" 11 11, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313b170 .functor NAND 1, L_0x5c7c3313b6c0, L_0x5c7c3313b7b0, C4<1>, C4<1>;
v0x5c7c32f0f240_0 .net "in_a", 0 0, L_0x5c7c3313b6c0;  1 drivers
v0x5c7c32f0f320_0 .net "in_b", 0 0, L_0x5c7c3313b7b0;  1 drivers
v0x5c7c32f0f3e0_0 .net "out", 0 0, L_0x5c7c3313b170;  1 drivers
S_0x5c7c32f0f530 .scope module, "nand_gate8" "Nand" 11 12, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313b930 .functor NAND 1, L_0x5c7c3313b9a0, L_0x5c7c3313ba90, C4<1>, C4<1>;
v0x5c7c32f0f760_0 .net "in_a", 0 0, L_0x5c7c3313b9a0;  1 drivers
v0x5c7c32f0f840_0 .net "in_b", 0 0, L_0x5c7c3313ba90;  1 drivers
v0x5c7c32f0f900_0 .net "out", 0 0, L_0x5c7c3313b930;  1 drivers
S_0x5c7c32f0fa50 .scope module, "nand_gate9" "Nand" 11 13, 6 1 0, S_0x5c7c32f0aa20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313bc20 .functor NAND 1, L_0x5c7c3313bc90, L_0x5c7c3313bd80, C4<1>, C4<1>;
v0x5c7c32f0fc80_0 .net "in_a", 0 0, L_0x5c7c3313bc90;  1 drivers
v0x5c7c32f0fd60_0 .net "in_b", 0 0, L_0x5c7c3313bd80;  1 drivers
v0x5c7c32f0fe20_0 .net "out", 0 0, L_0x5c7c3313bc20;  1 drivers
S_0x5c7c32cd69b0 .scope module, "DMux4Way" "DMux4Way" 12 3;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in";
    .port_info 1 /INPUT 2 "sel";
    .port_info 2 /OUTPUT 1 "a";
    .port_info 3 /OUTPUT 1 "b";
    .port_info 4 /OUTPUT 1 "c";
    .port_info 5 /OUTPUT 1 "d";
v0x5c7c32f1b0e0_0 .net "a", 0 0, L_0x5c7c3313db70;  1 drivers
v0x5c7c32f1b230_0 .net "b", 0 0, L_0x5c7c32f171b0;  1 drivers
v0x5c7c32f1b380_0 .net "c", 0 0, L_0x5c7c3313de20;  1 drivers
v0x5c7c32f1b4b0_0 .net "d", 0 0, L_0x5c7c32f1aac0;  1 drivers
o0x7d2eeb862198 .functor BUFZ 1, C4<z>; HiZ drive
v0x5c7c32f1b5e0_0 .net "in", 0 0, o0x7d2eeb862198;  0 drivers
o0x7d2eeb863698 .functor BUFZ 2, C4<zz>; HiZ drive
v0x5c7c32f1b680_0 .net "sel", 1 0, o0x7d2eeb863698;  0 drivers
v0x5c7c32f1b720_0 .net "tmp_ab", 0 0, L_0x5c7c3313d8a0;  1 drivers
v0x5c7c32f1b7c0_0 .net "tmp_cd", 0 0, L_0x5c7c3313d980;  1 drivers
L_0x5c7c3313d9f0 .part o0x7d2eeb863698, 1, 1;
L_0x5c7c3313dc50 .part o0x7d2eeb863698, 0, 1;
L_0x5c7c3313e010 .part o0x7d2eeb863698, 0, 1;
S_0x5c7c32f10580 .scope module, "dmux_gate1" "DMux" 12 7, 13 2 0, S_0x5c7c32cd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in";
    .port_info 1 /OUTPUT 1 "out_a";
    .port_info 2 /OUTPUT 1 "out_b";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f13a80_0 .net "in", 0 0, o0x7d2eeb862198;  alias, 0 drivers
v0x5c7c32f13bb0_0 .net "out_a", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f13c70_0 .net "out_b", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f13d10_0 .net "sel", 0 0, L_0x5c7c3313d9f0;  1 drivers
v0x5c7c32f13db0_0 .net "sel_out", 0 0, L_0x5c7c3313d7c0;  1 drivers
S_0x5c7c32f10800 .scope module, "and_gate" "And" 13 8, 5 2 0, S_0x5c7c32f10580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f118f0_0 .net "in_a", 0 0, o0x7d2eeb862198;  alias, 0 drivers
v0x5c7c32f119c0_0 .net "in_b", 0 0, L_0x5c7c3313d7c0;  alias, 1 drivers
v0x5c7c32f11a90_0 .net "out", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f11bb0_0 .net "temp_out", 0 0, L_0x5c7c3313d830;  1 drivers
S_0x5c7c32f10a70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f10800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313d830 .functor NAND 1, o0x7d2eeb862198, L_0x5c7c3313d7c0, C4<1>, C4<1>;
v0x5c7c32f10ce0_0 .net "in_a", 0 0, o0x7d2eeb862198;  alias, 0 drivers
v0x5c7c32f10dc0_0 .net "in_b", 0 0, L_0x5c7c3313d7c0;  alias, 1 drivers
v0x5c7c32f10e80_0 .net "out", 0 0, L_0x5c7c3313d830;  alias, 1 drivers
S_0x5c7c32f10fd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f10800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f11740_0 .net "in_a", 0 0, L_0x5c7c3313d830;  alias, 1 drivers
v0x5c7c32f117e0_0 .net "out", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
S_0x5c7c32f111f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f10fd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313d8a0 .functor NAND 1, L_0x5c7c3313d830, L_0x5c7c3313d830, C4<1>, C4<1>;
v0x5c7c32f11460_0 .net "in_a", 0 0, L_0x5c7c3313d830;  alias, 1 drivers
v0x5c7c32f11550_0 .net "in_b", 0 0, L_0x5c7c3313d830;  alias, 1 drivers
v0x5c7c32f11640_0 .net "out", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
S_0x5c7c32f11d00 .scope module, "and_gate3" "And" 13 9, 5 2 0, S_0x5c7c32f10580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f12d30_0 .net "in_a", 0 0, o0x7d2eeb862198;  alias, 0 drivers
v0x5c7c32f12dd0_0 .net "in_b", 0 0, L_0x5c7c3313d9f0;  alias, 1 drivers
v0x5c7c32f12ec0_0 .net "out", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f12fe0_0 .net "temp_out", 0 0, L_0x5c7c3313d910;  1 drivers
S_0x5c7c32f11ee0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f11d00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313d910 .functor NAND 1, o0x7d2eeb862198, L_0x5c7c3313d9f0, C4<1>, C4<1>;
v0x5c7c32f12150_0 .net "in_a", 0 0, o0x7d2eeb862198;  alias, 0 drivers
v0x5c7c32f12260_0 .net "in_b", 0 0, L_0x5c7c3313d9f0;  alias, 1 drivers
v0x5c7c32f12320_0 .net "out", 0 0, L_0x5c7c3313d910;  alias, 1 drivers
S_0x5c7c32f12440 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f11d00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f12b80_0 .net "in_a", 0 0, L_0x5c7c3313d910;  alias, 1 drivers
v0x5c7c32f12c20_0 .net "out", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
S_0x5c7c32f12660 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f12440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313d980 .functor NAND 1, L_0x5c7c3313d910, L_0x5c7c3313d910, C4<1>, C4<1>;
v0x5c7c32f128d0_0 .net "in_a", 0 0, L_0x5c7c3313d910;  alias, 1 drivers
v0x5c7c32f12990_0 .net "in_b", 0 0, L_0x5c7c3313d910;  alias, 1 drivers
v0x5c7c32f12a80_0 .net "out", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
S_0x5c7c32f13130 .scope module, "not_gate2" "Not" 13 7, 7 3 0, S_0x5c7c32f10580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f13850_0 .net "in_a", 0 0, L_0x5c7c3313d9f0;  alias, 1 drivers
v0x5c7c32f13980_0 .net "out", 0 0, L_0x5c7c3313d7c0;  alias, 1 drivers
S_0x5c7c32f13300 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f13130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313d7c0 .functor NAND 1, L_0x5c7c3313d9f0, L_0x5c7c3313d9f0, C4<1>, C4<1>;
v0x5c7c32f13550_0 .net "in_a", 0 0, L_0x5c7c3313d9f0;  alias, 1 drivers
v0x5c7c32f13660_0 .net "in_b", 0 0, L_0x5c7c3313d9f0;  alias, 1 drivers
v0x5c7c32f13720_0 .net "out", 0 0, L_0x5c7c3313d7c0;  alias, 1 drivers
S_0x5c7c32f13f20 .scope module, "dmux_gate2" "DMux" 12 8, 13 2 0, S_0x5c7c32cd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in";
    .port_info 1 /OUTPUT 1 "out_a";
    .port_info 2 /OUTPUT 1 "out_b";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f17340_0 .net "in", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f174f0_0 .net "out_a", 0 0, L_0x5c7c3313db70;  alias, 1 drivers
v0x5c7c32f175b0_0 .net "out_b", 0 0, L_0x5c7c32f171b0;  alias, 1 drivers
v0x5c7c32f17650_0 .net "sel", 0 0, L_0x5c7c3313dc50;  1 drivers
v0x5c7c32f176f0_0 .net "sel_out", 0 0, L_0x5c7c3313da90;  1 drivers
S_0x5c7c32f14140 .scope module, "and_gate" "And" 13 8, 5 2 0, S_0x5c7c32f13f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f151e0_0 .net "in_a", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f15280_0 .net "in_b", 0 0, L_0x5c7c3313da90;  alias, 1 drivers
v0x5c7c32f15370_0 .net "out", 0 0, L_0x5c7c3313db70;  alias, 1 drivers
v0x5c7c32f15490_0 .net "temp_out", 0 0, L_0x5c7c3313db00;  1 drivers
S_0x5c7c32f14340 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f14140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313db00 .functor NAND 1, L_0x5c7c3313d8a0, L_0x5c7c3313da90, C4<1>, C4<1>;
v0x5c7c32f145b0_0 .net "in_a", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f14700_0 .net "in_b", 0 0, L_0x5c7c3313da90;  alias, 1 drivers
v0x5c7c32f147c0_0 .net "out", 0 0, L_0x5c7c3313db00;  alias, 1 drivers
S_0x5c7c32f14910 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f14140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f15030_0 .net "in_a", 0 0, L_0x5c7c3313db00;  alias, 1 drivers
v0x5c7c32f150d0_0 .net "out", 0 0, L_0x5c7c3313db70;  alias, 1 drivers
S_0x5c7c32f14ae0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f14910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313db70 .functor NAND 1, L_0x5c7c3313db00, L_0x5c7c3313db00, C4<1>, C4<1>;
v0x5c7c32f14d50_0 .net "in_a", 0 0, L_0x5c7c3313db00;  alias, 1 drivers
v0x5c7c32f14e40_0 .net "in_b", 0 0, L_0x5c7c3313db00;  alias, 1 drivers
v0x5c7c32f14f30_0 .net "out", 0 0, L_0x5c7c3313db70;  alias, 1 drivers
S_0x5c7c32f155e0 .scope module, "and_gate3" "And" 13 9, 5 2 0, S_0x5c7c32f13f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f165f0_0 .net "in_a", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f16690_0 .net "in_b", 0 0, L_0x5c7c3313dc50;  alias, 1 drivers
v0x5c7c32f16780_0 .net "out", 0 0, L_0x5c7c32f171b0;  alias, 1 drivers
v0x5c7c32f168a0_0 .net "temp_out", 0 0, L_0x5c7c3313dbe0;  1 drivers
S_0x5c7c32f157c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f155e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313dbe0 .functor NAND 1, L_0x5c7c3313d8a0, L_0x5c7c3313dc50, C4<1>, C4<1>;
v0x5c7c32f15a30_0 .net "in_a", 0 0, L_0x5c7c3313d8a0;  alias, 1 drivers
v0x5c7c32f15af0_0 .net "in_b", 0 0, L_0x5c7c3313dc50;  alias, 1 drivers
v0x5c7c32f15bb0_0 .net "out", 0 0, L_0x5c7c3313dbe0;  alias, 1 drivers
S_0x5c7c32f15cd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f155e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f16440_0 .net "in_a", 0 0, L_0x5c7c3313dbe0;  alias, 1 drivers
v0x5c7c32f164e0_0 .net "out", 0 0, L_0x5c7c32f171b0;  alias, 1 drivers
S_0x5c7c32f15ef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f15cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f171b0 .functor NAND 1, L_0x5c7c3313dbe0, L_0x5c7c3313dbe0, C4<1>, C4<1>;
v0x5c7c32f16160_0 .net "in_a", 0 0, L_0x5c7c3313dbe0;  alias, 1 drivers
v0x5c7c32f16250_0 .net "in_b", 0 0, L_0x5c7c3313dbe0;  alias, 1 drivers
v0x5c7c32f16340_0 .net "out", 0 0, L_0x5c7c32f171b0;  alias, 1 drivers
S_0x5c7c32f169f0 .scope module, "not_gate2" "Not" 13 7, 7 3 0, S_0x5c7c32f13f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f17110_0 .net "in_a", 0 0, L_0x5c7c3313dc50;  alias, 1 drivers
v0x5c7c32f17240_0 .net "out", 0 0, L_0x5c7c3313da90;  alias, 1 drivers
S_0x5c7c32f16bc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f169f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313da90 .functor NAND 1, L_0x5c7c3313dc50, L_0x5c7c3313dc50, C4<1>, C4<1>;
v0x5c7c32f16e10_0 .net "in_a", 0 0, L_0x5c7c3313dc50;  alias, 1 drivers
v0x5c7c32f16f20_0 .net "in_b", 0 0, L_0x5c7c3313dc50;  alias, 1 drivers
v0x5c7c32f16fe0_0 .net "out", 0 0, L_0x5c7c3313da90;  alias, 1 drivers
S_0x5c7c32f177d0 .scope module, "dmux_gate3" "DMux" 12 9, 13 2 0, S_0x5c7c32cd69b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in";
    .port_info 1 /OUTPUT 1 "out_a";
    .port_info 2 /OUTPUT 1 "out_b";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f1ac50_0 .net "in", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f1ae00_0 .net "out_a", 0 0, L_0x5c7c3313de20;  alias, 1 drivers
v0x5c7c32f1aec0_0 .net "out_b", 0 0, L_0x5c7c32f1aac0;  alias, 1 drivers
v0x5c7c32f1af60_0 .net "sel", 0 0, L_0x5c7c3313e010;  1 drivers
v0x5c7c32f1b000_0 .net "sel_out", 0 0, L_0x5c7c3313dd40;  1 drivers
S_0x5c7c32f17a00 .scope module, "and_gate" "And" 13 8, 5 2 0, S_0x5c7c32f177d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f18af0_0 .net "in_a", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f18b90_0 .net "in_b", 0 0, L_0x5c7c3313dd40;  alias, 1 drivers
v0x5c7c32f18c80_0 .net "out", 0 0, L_0x5c7c3313de20;  alias, 1 drivers
v0x5c7c32f18da0_0 .net "temp_out", 0 0, L_0x5c7c3313ddb0;  1 drivers
S_0x5c7c32f17c50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f17a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313ddb0 .functor NAND 1, L_0x5c7c3313d980, L_0x5c7c3313dd40, C4<1>, C4<1>;
v0x5c7c32f17ec0_0 .net "in_a", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f18010_0 .net "in_b", 0 0, L_0x5c7c3313dd40;  alias, 1 drivers
v0x5c7c32f180d0_0 .net "out", 0 0, L_0x5c7c3313ddb0;  alias, 1 drivers
S_0x5c7c32f18220 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f17a00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f18940_0 .net "in_a", 0 0, L_0x5c7c3313ddb0;  alias, 1 drivers
v0x5c7c32f189e0_0 .net "out", 0 0, L_0x5c7c3313de20;  alias, 1 drivers
S_0x5c7c32f183f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f18220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313de20 .functor NAND 1, L_0x5c7c3313ddb0, L_0x5c7c3313ddb0, C4<1>, C4<1>;
v0x5c7c32f18660_0 .net "in_a", 0 0, L_0x5c7c3313ddb0;  alias, 1 drivers
v0x5c7c32f18750_0 .net "in_b", 0 0, L_0x5c7c3313ddb0;  alias, 1 drivers
v0x5c7c32f18840_0 .net "out", 0 0, L_0x5c7c3313de20;  alias, 1 drivers
S_0x5c7c32f18ef0 .scope module, "and_gate3" "And" 13 9, 5 2 0, S_0x5c7c32f177d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f19f00_0 .net "in_a", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f19fa0_0 .net "in_b", 0 0, L_0x5c7c3313e010;  alias, 1 drivers
v0x5c7c32f1a090_0 .net "out", 0 0, L_0x5c7c32f1aac0;  alias, 1 drivers
v0x5c7c32f1a1b0_0 .net "temp_out", 0 0, L_0x5c7c3313de90;  1 drivers
S_0x5c7c32f190d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f18ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313de90 .functor NAND 1, L_0x5c7c3313d980, L_0x5c7c3313e010, C4<1>, C4<1>;
v0x5c7c32f19340_0 .net "in_a", 0 0, L_0x5c7c3313d980;  alias, 1 drivers
v0x5c7c32f19400_0 .net "in_b", 0 0, L_0x5c7c3313e010;  alias, 1 drivers
v0x5c7c32f194c0_0 .net "out", 0 0, L_0x5c7c3313de90;  alias, 1 drivers
S_0x5c7c32f195e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f18ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f19d50_0 .net "in_a", 0 0, L_0x5c7c3313de90;  alias, 1 drivers
v0x5c7c32f19df0_0 .net "out", 0 0, L_0x5c7c32f1aac0;  alias, 1 drivers
S_0x5c7c32f19800 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f195e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f1aac0 .functor NAND 1, L_0x5c7c3313de90, L_0x5c7c3313de90, C4<1>, C4<1>;
v0x5c7c32f19a70_0 .net "in_a", 0 0, L_0x5c7c3313de90;  alias, 1 drivers
v0x5c7c32f19b60_0 .net "in_b", 0 0, L_0x5c7c3313de90;  alias, 1 drivers
v0x5c7c32f19c50_0 .net "out", 0 0, L_0x5c7c32f1aac0;  alias, 1 drivers
S_0x5c7c32f1a300 .scope module, "not_gate2" "Not" 13 7, 7 3 0, S_0x5c7c32f177d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f1aa20_0 .net "in_a", 0 0, L_0x5c7c3313e010;  alias, 1 drivers
v0x5c7c32f1ab50_0 .net "out", 0 0, L_0x5c7c3313dd40;  alias, 1 drivers
S_0x5c7c32f1a4d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f1a300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313dd40 .functor NAND 1, L_0x5c7c3313e010, L_0x5c7c3313e010, C4<1>, C4<1>;
v0x5c7c32f1a720_0 .net "in_a", 0 0, L_0x5c7c3313e010;  alias, 1 drivers
v0x5c7c32f1a830_0 .net "in_b", 0 0, L_0x5c7c3313e010;  alias, 1 drivers
v0x5c7c32f1a8f0_0 .net "out", 0 0, L_0x5c7c3313dd40;  alias, 1 drivers
S_0x5c7c32cac1f0 .scope module, "Mux4Way16" "Mux4Way16" 14 3;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "in_a";
    .port_info 1 /INPUT 16 "in_b";
    .port_info 2 /INPUT 16 "in_c";
    .port_info 3 /INPUT 16 "in_d";
    .port_info 4 /OUTPUT 16 "out";
    .port_info 5 /INPUT 2 "sel";
v0x5c7c33111490_0 .net "group_1", 15 0, L_0x5c7c3314c880;  1 drivers
v0x5c7c331115c0_0 .net "group_2", 15 0, L_0x5c7c3315b4e0;  1 drivers
o0x7d2eeb875e18 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c331116d0_0 .net "in_a", 15 0, o0x7d2eeb875e18;  0 drivers
o0x7d2eeb8885c8 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c33111770_0 .net "in_b", 15 0, o0x7d2eeb8885c8;  0 drivers
o0x7d2eeb875e48 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c33111810_0 .net "in_c", 15 0, o0x7d2eeb875e48;  0 drivers
o0x7d2eeb8885f8 .functor BUFZ 16, C4<zzzzzzzzzzzzzzzz>; HiZ drive
v0x5c7c33111900_0 .net "in_d", 15 0, o0x7d2eeb8885f8;  0 drivers
v0x5c7c331119a0_0 .net "out", 15 0, L_0x5c7c33169f80;  1 drivers
o0x7d2eeb839e98 .functor BUFZ 2, C4<zz>; HiZ drive
v0x5c7c33111a70_0 .net "sel", 1 0, o0x7d2eeb839e98;  0 drivers
L_0x5c7c3314c910 .part o0x7d2eeb839e98, 1, 1;
L_0x5c7c3315b570 .part o0x7d2eeb839e98, 1, 1;
L_0x5c7c33169ff0 .part o0x7d2eeb839e98, 0, 1;
S_0x5c7c32f1b960 .scope module, "mux16_gate1" "Mux16" 14 13, 15 3 0, S_0x5c7c32cac1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "in_a";
    .port_info 1 /INPUT 16 "in_b";
    .port_info 2 /OUTPUT 16 "out";
    .port_info 3 /INPUT 1 "sel";
L_0x5c7c3314c880 .functor BUFZ 16, L_0x5c7c3314c7e0, C4<0000000000000000>, C4<0000000000000000>, C4<0000000000000000>;
v0x5c7c32fb8240_0 .net "in_a", 15 0, o0x7d2eeb875e18;  alias, 0 drivers
v0x5c7c32fb8340_0 .net "in_b", 15 0, o0x7d2eeb875e48;  alias, 0 drivers
v0x5c7c32fb8420_0 .net "out", 15 0, L_0x5c7c3314c880;  alias, 1 drivers
v0x5c7c32fb84e0_0 .net "sel", 0 0, L_0x5c7c3314c910;  1 drivers
v0x5c7c32fb8580_0 .net/s "tmp_out", 15 0, L_0x5c7c3314c7e0;  1 drivers
L_0x5c7c3313eb80 .part o0x7d2eeb875e18, 0, 1;
L_0x5c7c3313ec40 .part o0x7d2eeb875e48, 0, 1;
L_0x5c7c3313f9b0 .part o0x7d2eeb875e18, 1, 1;
L_0x5c7c3313fa50 .part o0x7d2eeb875e48, 1, 1;
L_0x5c7c331407a0 .part o0x7d2eeb875e18, 2, 1;
L_0x5c7c33140840 .part o0x7d2eeb875e48, 2, 1;
L_0x5c7c331415f0 .part o0x7d2eeb875e18, 3, 1;
L_0x5c7c33141690 .part o0x7d2eeb875e48, 3, 1;
L_0x5c7c33142400 .part o0x7d2eeb875e18, 4, 1;
L_0x5c7c331424a0 .part o0x7d2eeb875e48, 4, 1;
L_0x5c7c33143270 .part o0x7d2eeb875e18, 5, 1;
L_0x5c7c33143310 .part o0x7d2eeb875e48, 5, 1;
L_0x5c7c331440f0 .part o0x7d2eeb875e18, 6, 1;
L_0x5c7c331442a0 .part o0x7d2eeb875e48, 6, 1;
L_0x5c7c33145130 .part o0x7d2eeb875e18, 7, 1;
L_0x5c7c331451d0 .part o0x7d2eeb875e48, 7, 1;
L_0x5c7c33145fd0 .part o0x7d2eeb875e18, 8, 1;
L_0x5c7c33146070 .part o0x7d2eeb875e48, 8, 1;
L_0x5c7c33146df0 .part o0x7d2eeb875e18, 9, 1;
L_0x5c7c33146e90 .part o0x7d2eeb875e48, 9, 1;
L_0x5c7c33146110 .part o0x7d2eeb875e18, 10, 1;
L_0x5c7c331483f0 .part o0x7d2eeb875e48, 10, 1;
L_0x5c7c33148ea0 .part o0x7d2eeb875e18, 11, 1;
L_0x5c7c33148f40 .part o0x7d2eeb875e48, 11, 1;
L_0x5c7c33149a00 .part o0x7d2eeb875e18, 12, 1;
L_0x5c7c33149aa0 .part o0x7d2eeb875e48, 12, 1;
L_0x5c7c3314a790 .part o0x7d2eeb875e18, 13, 1;
L_0x5c7c3314a830 .part o0x7d2eeb875e48, 13, 1;
L_0x5c7c3314b690 .part o0x7d2eeb875e18, 14, 1;
L_0x5c7c3314b730 .part o0x7d2eeb875e48, 14, 1;
L_0x5c7c3314c590 .part o0x7d2eeb875e18, 15, 1;
L_0x5c7c3314c630 .part o0x7d2eeb875e48, 15, 1;
LS_0x5c7c3314c7e0_0_0 .concat8 [ 1 1 1 1], L_0x5c7c3313e9c0, L_0x5c7c3313f7f0, L_0x5c7c331405e0, L_0x5c7c33141430;
LS_0x5c7c3314c7e0_0_4 .concat8 [ 1 1 1 1], L_0x5c7c33142240, L_0x5c7c331430b0, L_0x5c7c33143f30, L_0x5c7c33144f70;
LS_0x5c7c3314c7e0_0_8 .concat8 [ 1 1 1 1], L_0x5c7c33145e10, L_0x5c7c33146c30, L_0x5c7c33148270, L_0x5c7c33148d20;
LS_0x5c7c3314c7e0_0_12 .concat8 [ 1 1 1 1], L_0x5c7c33149880, L_0x5c7c3314a5d0, L_0x5c7c3314b4d0, L_0x5c7c3314c3d0;
L_0x5c7c3314c7e0 .concat8 [ 4 4 4 4], LS_0x5c7c3314c7e0_0_0, LS_0x5c7c3314c7e0_0_4, LS_0x5c7c3314c7e0_0_8, LS_0x5c7c3314c7e0_0_12;
S_0x5c7c32f1bb80 .scope module, "mux_gate0" "Mux" 15 7, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f25090_0 .net "in_a", 0 0, L_0x5c7c3313eb80;  1 drivers
v0x5c7c32f25130_0 .net "in_b", 0 0, L_0x5c7c3313ec40;  1 drivers
v0x5c7c32f25240_0 .net "out", 0 0, L_0x5c7c3313e9c0;  1 drivers
v0x5c7c32f252e0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f25380_0 .net "sel_out", 0 0, L_0x5c7c3313e0b0;  1 drivers
v0x5c7c32f25500_0 .net "temp_a_out", 0 0, L_0x5c7c3313e190;  1 drivers
v0x5c7c32f256b0_0 .net "temp_b_out", 0 0, L_0x5c7c3313e290;  1 drivers
S_0x5c7c32f1bdd0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f1bb80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f1cde0_0 .net "in_a", 0 0, L_0x5c7c3313eb80;  alias, 1 drivers
v0x5c7c32f1ceb0_0 .net "in_b", 0 0, L_0x5c7c3313e0b0;  alias, 1 drivers
v0x5c7c32f1cf80_0 .net "out", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
v0x5c7c32f1d0a0_0 .net "temp_out", 0 0, L_0x5c7c3313e120;  1 drivers
S_0x5c7c32f1bfa0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f1bdd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e120 .functor NAND 1, L_0x5c7c3313eb80, L_0x5c7c3313e0b0, C4<1>, C4<1>;
v0x5c7c32f1c210_0 .net "in_a", 0 0, L_0x5c7c3313eb80;  alias, 1 drivers
v0x5c7c32f1c2f0_0 .net "in_b", 0 0, L_0x5c7c3313e0b0;  alias, 1 drivers
v0x5c7c32f1c3b0_0 .net "out", 0 0, L_0x5c7c3313e120;  alias, 1 drivers
S_0x5c7c32f1c500 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f1bdd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f1cc30_0 .net "in_a", 0 0, L_0x5c7c3313e120;  alias, 1 drivers
v0x5c7c32f1ccd0_0 .net "out", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
S_0x5c7c32f1c6e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f1c500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e190 .functor NAND 1, L_0x5c7c3313e120, L_0x5c7c3313e120, C4<1>, C4<1>;
v0x5c7c32f1c950_0 .net "in_a", 0 0, L_0x5c7c3313e120;  alias, 1 drivers
v0x5c7c32f1ca40_0 .net "in_b", 0 0, L_0x5c7c3313e120;  alias, 1 drivers
v0x5c7c32f1cb30_0 .net "out", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
S_0x5c7c32f1d1f0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f1bb80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f1e220_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f1e2f0_0 .net "in_b", 0 0, L_0x5c7c3313ec40;  alias, 1 drivers
v0x5c7c32f1e3c0_0 .net "out", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
v0x5c7c32f1e4e0_0 .net "temp_out", 0 0, L_0x5c7c3313e200;  1 drivers
S_0x5c7c32f1d3d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f1d1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e200 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3313ec40, C4<1>, C4<1>;
v0x5c7c32f1d640_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f1d720_0 .net "in_b", 0 0, L_0x5c7c3313ec40;  alias, 1 drivers
v0x5c7c32f1d7e0_0 .net "out", 0 0, L_0x5c7c3313e200;  alias, 1 drivers
S_0x5c7c32f1d900 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f1d1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f1e070_0 .net "in_a", 0 0, L_0x5c7c3313e200;  alias, 1 drivers
v0x5c7c32f1e110_0 .net "out", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
S_0x5c7c32f1db20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f1d900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e290 .functor NAND 1, L_0x5c7c3313e200, L_0x5c7c3313e200, C4<1>, C4<1>;
v0x5c7c32f1dd90_0 .net "in_a", 0 0, L_0x5c7c3313e200;  alias, 1 drivers
v0x5c7c32f1de80_0 .net "in_b", 0 0, L_0x5c7c3313e200;  alias, 1 drivers
v0x5c7c32f1df70_0 .net "out", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
S_0x5c7c32f1e630 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f1bb80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f1ed50_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f1ee80_0 .net "out", 0 0, L_0x5c7c3313e0b0;  alias, 1 drivers
S_0x5c7c32f1e800 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f1e630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e0b0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f1ea50_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f1eb60_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f1ec20_0 .net "out", 0 0, L_0x5c7c3313e0b0;  alias, 1 drivers
S_0x5c7c32f1ef80 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f1bb80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f249e0_0 .net "branch1_out", 0 0, L_0x5c7c3313e4a0;  1 drivers
v0x5c7c32f24b10_0 .net "branch2_out", 0 0, L_0x5c7c3313e730;  1 drivers
v0x5c7c32f24c60_0 .net "in_a", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
v0x5c7c32f24d30_0 .net "in_b", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
v0x5c7c32f24dd0_0 .net "out", 0 0, L_0x5c7c3313e9c0;  alias, 1 drivers
v0x5c7c32f24e70_0 .net "temp1_out", 0 0, L_0x5c7c3313e3f0;  1 drivers
v0x5c7c32f24f10_0 .net "temp2_out", 0 0, L_0x5c7c3313e680;  1 drivers
v0x5c7c32f24fb0_0 .net "temp3_out", 0 0, L_0x5c7c3313e910;  1 drivers
S_0x5c7c32f1f160 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f1ef80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f20220_0 .net "in_a", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
v0x5c7c32f202c0_0 .net "in_b", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
v0x5c7c32f20380_0 .net "out", 0 0, L_0x5c7c3313e3f0;  alias, 1 drivers
v0x5c7c32f204a0_0 .net "temp_out", 0 0, L_0x5c7c3313e340;  1 drivers
S_0x5c7c32f1f3d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f1f160;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e340 .functor NAND 1, L_0x5c7c3313e190, L_0x5c7c3313e190, C4<1>, C4<1>;
v0x5c7c32f1f640_0 .net "in_a", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
v0x5c7c32f1f700_0 .net "in_b", 0 0, L_0x5c7c3313e190;  alias, 1 drivers
v0x5c7c32f1f850_0 .net "out", 0 0, L_0x5c7c3313e340;  alias, 1 drivers
S_0x5c7c32f1f950 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f1f160;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f20070_0 .net "in_a", 0 0, L_0x5c7c3313e340;  alias, 1 drivers
v0x5c7c32f20110_0 .net "out", 0 0, L_0x5c7c3313e3f0;  alias, 1 drivers
S_0x5c7c32f1fb20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f1f950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e3f0 .functor NAND 1, L_0x5c7c3313e340, L_0x5c7c3313e340, C4<1>, C4<1>;
v0x5c7c32f1fd90_0 .net "in_a", 0 0, L_0x5c7c3313e340;  alias, 1 drivers
v0x5c7c32f1fe80_0 .net "in_b", 0 0, L_0x5c7c3313e340;  alias, 1 drivers
v0x5c7c32f1ff70_0 .net "out", 0 0, L_0x5c7c3313e3f0;  alias, 1 drivers
S_0x5c7c32f20610 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f1ef80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f21640_0 .net "in_a", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
v0x5c7c32f216e0_0 .net "in_b", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
v0x5c7c32f217a0_0 .net "out", 0 0, L_0x5c7c3313e680;  alias, 1 drivers
v0x5c7c32f218c0_0 .net "temp_out", 0 0, L_0x5c7c32f23460;  1 drivers
S_0x5c7c32f207f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f20610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f23460 .functor NAND 1, L_0x5c7c3313e290, L_0x5c7c3313e290, C4<1>, C4<1>;
v0x5c7c32f20a60_0 .net "in_a", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
v0x5c7c32f20b20_0 .net "in_b", 0 0, L_0x5c7c3313e290;  alias, 1 drivers
v0x5c7c32f20c70_0 .net "out", 0 0, L_0x5c7c32f23460;  alias, 1 drivers
S_0x5c7c32f20d70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f20610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f21490_0 .net "in_a", 0 0, L_0x5c7c32f23460;  alias, 1 drivers
v0x5c7c32f21530_0 .net "out", 0 0, L_0x5c7c3313e680;  alias, 1 drivers
S_0x5c7c32f20f40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f20d70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e680 .functor NAND 1, L_0x5c7c32f23460, L_0x5c7c32f23460, C4<1>, C4<1>;
v0x5c7c32f211b0_0 .net "in_a", 0 0, L_0x5c7c32f23460;  alias, 1 drivers
v0x5c7c32f212a0_0 .net "in_b", 0 0, L_0x5c7c32f23460;  alias, 1 drivers
v0x5c7c32f21390_0 .net "out", 0 0, L_0x5c7c3313e680;  alias, 1 drivers
S_0x5c7c32f21a30 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f1ef80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f22a70_0 .net "in_a", 0 0, L_0x5c7c3313e4a0;  alias, 1 drivers
v0x5c7c32f22b40_0 .net "in_b", 0 0, L_0x5c7c3313e730;  alias, 1 drivers
v0x5c7c32f22c10_0 .net "out", 0 0, L_0x5c7c3313e910;  alias, 1 drivers
v0x5c7c32f22d30_0 .net "temp_out", 0 0, L_0x5c7c32f23dd0;  1 drivers
S_0x5c7c32f21c10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f21a30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f23dd0 .functor NAND 1, L_0x5c7c3313e4a0, L_0x5c7c3313e730, C4<1>, C4<1>;
v0x5c7c32f21e60_0 .net "in_a", 0 0, L_0x5c7c3313e4a0;  alias, 1 drivers
v0x5c7c32f21f40_0 .net "in_b", 0 0, L_0x5c7c3313e730;  alias, 1 drivers
v0x5c7c32f22000_0 .net "out", 0 0, L_0x5c7c32f23dd0;  alias, 1 drivers
S_0x5c7c32f22150 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f21a30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f228c0_0 .net "in_a", 0 0, L_0x5c7c32f23dd0;  alias, 1 drivers
v0x5c7c32f22960_0 .net "out", 0 0, L_0x5c7c3313e910;  alias, 1 drivers
S_0x5c7c32f22370 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f22150;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e910 .functor NAND 1, L_0x5c7c32f23dd0, L_0x5c7c32f23dd0, C4<1>, C4<1>;
v0x5c7c32f225e0_0 .net "in_a", 0 0, L_0x5c7c32f23dd0;  alias, 1 drivers
v0x5c7c32f226d0_0 .net "in_b", 0 0, L_0x5c7c32f23dd0;  alias, 1 drivers
v0x5c7c32f227c0_0 .net "out", 0 0, L_0x5c7c3313e910;  alias, 1 drivers
S_0x5c7c32f22e80 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f1ef80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f235b0_0 .net "in_a", 0 0, L_0x5c7c3313e3f0;  alias, 1 drivers
v0x5c7c32f23650_0 .net "out", 0 0, L_0x5c7c3313e4a0;  alias, 1 drivers
S_0x5c7c32f23050 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f22e80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e4a0 .functor NAND 1, L_0x5c7c3313e3f0, L_0x5c7c3313e3f0, C4<1>, C4<1>;
v0x5c7c32f232c0_0 .net "in_a", 0 0, L_0x5c7c3313e3f0;  alias, 1 drivers
v0x5c7c32f23380_0 .net "in_b", 0 0, L_0x5c7c3313e3f0;  alias, 1 drivers
v0x5c7c32f234d0_0 .net "out", 0 0, L_0x5c7c3313e4a0;  alias, 1 drivers
S_0x5c7c32f23750 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f1ef80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f23f20_0 .net "in_a", 0 0, L_0x5c7c3313e680;  alias, 1 drivers
v0x5c7c32f23fc0_0 .net "out", 0 0, L_0x5c7c3313e730;  alias, 1 drivers
S_0x5c7c32f239c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f23750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e730 .functor NAND 1, L_0x5c7c3313e680, L_0x5c7c3313e680, C4<1>, C4<1>;
v0x5c7c32f23c30_0 .net "in_a", 0 0, L_0x5c7c3313e680;  alias, 1 drivers
v0x5c7c32f23cf0_0 .net "in_b", 0 0, L_0x5c7c3313e680;  alias, 1 drivers
v0x5c7c32f23e40_0 .net "out", 0 0, L_0x5c7c3313e730;  alias, 1 drivers
S_0x5c7c32f240c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f1ef80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f24860_0 .net "in_a", 0 0, L_0x5c7c3313e910;  alias, 1 drivers
v0x5c7c32f24900_0 .net "out", 0 0, L_0x5c7c3313e9c0;  alias, 1 drivers
S_0x5c7c32f242e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f240c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313e9c0 .functor NAND 1, L_0x5c7c3313e910, L_0x5c7c3313e910, C4<1>, C4<1>;
v0x5c7c32f24550_0 .net "in_a", 0 0, L_0x5c7c3313e910;  alias, 1 drivers
v0x5c7c32f24610_0 .net "in_b", 0 0, L_0x5c7c3313e910;  alias, 1 drivers
v0x5c7c32f24760_0 .net "out", 0 0, L_0x5c7c3313e9c0;  alias, 1 drivers
S_0x5c7c32f258a0 .scope module, "mux_gate1" "Mux" 15 8, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f2ec80_0 .net "in_a", 0 0, L_0x5c7c3313f9b0;  1 drivers
v0x5c7c32f2ed20_0 .net "in_b", 0 0, L_0x5c7c3313fa50;  1 drivers
v0x5c7c32f2ee30_0 .net "out", 0 0, L_0x5c7c3313f7f0;  1 drivers
v0x5c7c32f2eed0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f2ef70_0 .net "sel_out", 0 0, L_0x5c7c3313ece0;  1 drivers
v0x5c7c32f2f0f0_0 .net "temp_a_out", 0 0, L_0x5c7c3313ee40;  1 drivers
v0x5c7c32f2f2a0_0 .net "temp_b_out", 0 0, L_0x5c7c3313efa0;  1 drivers
S_0x5c7c32f25ac0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f258a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f26b00_0 .net "in_a", 0 0, L_0x5c7c3313f9b0;  alias, 1 drivers
v0x5c7c32f26bd0_0 .net "in_b", 0 0, L_0x5c7c3313ece0;  alias, 1 drivers
v0x5c7c32f26ca0_0 .net "out", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
v0x5c7c32f26dc0_0 .net "temp_out", 0 0, L_0x5c7c3313ed90;  1 drivers
S_0x5c7c32f25d10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f25ac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313ed90 .functor NAND 1, L_0x5c7c3313f9b0, L_0x5c7c3313ece0, C4<1>, C4<1>;
v0x5c7c32f25f80_0 .net "in_a", 0 0, L_0x5c7c3313f9b0;  alias, 1 drivers
v0x5c7c32f26060_0 .net "in_b", 0 0, L_0x5c7c3313ece0;  alias, 1 drivers
v0x5c7c32f26120_0 .net "out", 0 0, L_0x5c7c3313ed90;  alias, 1 drivers
S_0x5c7c32f26240 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f25ac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f26980_0 .net "in_a", 0 0, L_0x5c7c3313ed90;  alias, 1 drivers
v0x5c7c32f26a20_0 .net "out", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
S_0x5c7c32f26460 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f26240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313ee40 .functor NAND 1, L_0x5c7c3313ed90, L_0x5c7c3313ed90, C4<1>, C4<1>;
v0x5c7c32f266d0_0 .net "in_a", 0 0, L_0x5c7c3313ed90;  alias, 1 drivers
v0x5c7c32f26790_0 .net "in_b", 0 0, L_0x5c7c3313ed90;  alias, 1 drivers
v0x5c7c32f26880_0 .net "out", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
S_0x5c7c32f26e80 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f258a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f27e90_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f27f30_0 .net "in_b", 0 0, L_0x5c7c3313fa50;  alias, 1 drivers
v0x5c7c32f28020_0 .net "out", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
v0x5c7c32f28140_0 .net "temp_out", 0 0, L_0x5c7c3313eef0;  1 drivers
S_0x5c7c32f27060 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f26e80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313eef0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3313fa50, C4<1>, C4<1>;
v0x5c7c32f272d0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f27390_0 .net "in_b", 0 0, L_0x5c7c3313fa50;  alias, 1 drivers
v0x5c7c32f27450_0 .net "out", 0 0, L_0x5c7c3313eef0;  alias, 1 drivers
S_0x5c7c32f27570 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f26e80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f27ce0_0 .net "in_a", 0 0, L_0x5c7c3313eef0;  alias, 1 drivers
v0x5c7c32f27d80_0 .net "out", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
S_0x5c7c32f27790 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f27570;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313efa0 .functor NAND 1, L_0x5c7c3313eef0, L_0x5c7c3313eef0, C4<1>, C4<1>;
v0x5c7c32f27a00_0 .net "in_a", 0 0, L_0x5c7c3313eef0;  alias, 1 drivers
v0x5c7c32f27af0_0 .net "in_b", 0 0, L_0x5c7c3313eef0;  alias, 1 drivers
v0x5c7c32f27be0_0 .net "out", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
S_0x5c7c32f28200 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f258a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f28a10_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f28ab0_0 .net "out", 0 0, L_0x5c7c3313ece0;  alias, 1 drivers
S_0x5c7c32f283d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f28200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313ece0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f28620_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f287f0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f288b0_0 .net "out", 0 0, L_0x5c7c3313ece0;  alias, 1 drivers
S_0x5c7c32f28bb0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f258a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f2e5d0_0 .net "branch1_out", 0 0, L_0x5c7c3313f1b0;  1 drivers
v0x5c7c32f2e700_0 .net "branch2_out", 0 0, L_0x5c7c3313f4d0;  1 drivers
v0x5c7c32f2e850_0 .net "in_a", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
v0x5c7c32f2e920_0 .net "in_b", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
v0x5c7c32f2e9c0_0 .net "out", 0 0, L_0x5c7c3313f7f0;  alias, 1 drivers
v0x5c7c32f2ea60_0 .net "temp1_out", 0 0, L_0x5c7c3313f100;  1 drivers
v0x5c7c32f2eb00_0 .net "temp2_out", 0 0, L_0x5c7c3313f420;  1 drivers
v0x5c7c32f2eba0_0 .net "temp3_out", 0 0, L_0x5c7c3313f740;  1 drivers
S_0x5c7c32f28de0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f28bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f29e10_0 .net "in_a", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
v0x5c7c32f29eb0_0 .net "in_b", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
v0x5c7c32f29f70_0 .net "out", 0 0, L_0x5c7c3313f100;  alias, 1 drivers
v0x5c7c32f2a090_0 .net "temp_out", 0 0, L_0x5c7c3313f050;  1 drivers
S_0x5c7c32f29050 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f28de0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f050 .functor NAND 1, L_0x5c7c3313ee40, L_0x5c7c3313ee40, C4<1>, C4<1>;
v0x5c7c32f292c0_0 .net "in_a", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
v0x5c7c32f29380_0 .net "in_b", 0 0, L_0x5c7c3313ee40;  alias, 1 drivers
v0x5c7c32f29440_0 .net "out", 0 0, L_0x5c7c3313f050;  alias, 1 drivers
S_0x5c7c32f29540 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f28de0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f29c60_0 .net "in_a", 0 0, L_0x5c7c3313f050;  alias, 1 drivers
v0x5c7c32f29d00_0 .net "out", 0 0, L_0x5c7c3313f100;  alias, 1 drivers
S_0x5c7c32f29710 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f29540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f100 .functor NAND 1, L_0x5c7c3313f050, L_0x5c7c3313f050, C4<1>, C4<1>;
v0x5c7c32f29980_0 .net "in_a", 0 0, L_0x5c7c3313f050;  alias, 1 drivers
v0x5c7c32f29a70_0 .net "in_b", 0 0, L_0x5c7c3313f050;  alias, 1 drivers
v0x5c7c32f29b60_0 .net "out", 0 0, L_0x5c7c3313f100;  alias, 1 drivers
S_0x5c7c32f2a200 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f28bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f2b230_0 .net "in_a", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
v0x5c7c32f2b2d0_0 .net "in_b", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
v0x5c7c32f2b390_0 .net "out", 0 0, L_0x5c7c3313f420;  alias, 1 drivers
v0x5c7c32f2b4b0_0 .net "temp_out", 0 0, L_0x5c7c3313f370;  1 drivers
S_0x5c7c32f2a3e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f2a200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f370 .functor NAND 1, L_0x5c7c3313efa0, L_0x5c7c3313efa0, C4<1>, C4<1>;
v0x5c7c32f2a650_0 .net "in_a", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
v0x5c7c32f2a710_0 .net "in_b", 0 0, L_0x5c7c3313efa0;  alias, 1 drivers
v0x5c7c32f2a860_0 .net "out", 0 0, L_0x5c7c3313f370;  alias, 1 drivers
S_0x5c7c32f2a960 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f2a200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f2b080_0 .net "in_a", 0 0, L_0x5c7c3313f370;  alias, 1 drivers
v0x5c7c32f2b120_0 .net "out", 0 0, L_0x5c7c3313f420;  alias, 1 drivers
S_0x5c7c32f2ab30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f2a960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f420 .functor NAND 1, L_0x5c7c3313f370, L_0x5c7c3313f370, C4<1>, C4<1>;
v0x5c7c32f2ada0_0 .net "in_a", 0 0, L_0x5c7c3313f370;  alias, 1 drivers
v0x5c7c32f2ae90_0 .net "in_b", 0 0, L_0x5c7c3313f370;  alias, 1 drivers
v0x5c7c32f2af80_0 .net "out", 0 0, L_0x5c7c3313f420;  alias, 1 drivers
S_0x5c7c32f2b620 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f28bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f2c660_0 .net "in_a", 0 0, L_0x5c7c3313f1b0;  alias, 1 drivers
v0x5c7c32f2c730_0 .net "in_b", 0 0, L_0x5c7c3313f4d0;  alias, 1 drivers
v0x5c7c32f2c800_0 .net "out", 0 0, L_0x5c7c3313f740;  alias, 1 drivers
v0x5c7c32f2c920_0 .net "temp_out", 0 0, L_0x5c7c3313f690;  1 drivers
S_0x5c7c32f2b800 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f2b620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f690 .functor NAND 1, L_0x5c7c3313f1b0, L_0x5c7c3313f4d0, C4<1>, C4<1>;
v0x5c7c32f2ba50_0 .net "in_a", 0 0, L_0x5c7c3313f1b0;  alias, 1 drivers
v0x5c7c32f2bb30_0 .net "in_b", 0 0, L_0x5c7c3313f4d0;  alias, 1 drivers
v0x5c7c32f2bbf0_0 .net "out", 0 0, L_0x5c7c3313f690;  alias, 1 drivers
S_0x5c7c32f2bd40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f2b620;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f2c4b0_0 .net "in_a", 0 0, L_0x5c7c3313f690;  alias, 1 drivers
v0x5c7c32f2c550_0 .net "out", 0 0, L_0x5c7c3313f740;  alias, 1 drivers
S_0x5c7c32f2bf60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f2bd40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f740 .functor NAND 1, L_0x5c7c3313f690, L_0x5c7c3313f690, C4<1>, C4<1>;
v0x5c7c32f2c1d0_0 .net "in_a", 0 0, L_0x5c7c3313f690;  alias, 1 drivers
v0x5c7c32f2c2c0_0 .net "in_b", 0 0, L_0x5c7c3313f690;  alias, 1 drivers
v0x5c7c32f2c3b0_0 .net "out", 0 0, L_0x5c7c3313f740;  alias, 1 drivers
S_0x5c7c32f2ca70 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f28bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f2d1a0_0 .net "in_a", 0 0, L_0x5c7c3313f100;  alias, 1 drivers
v0x5c7c32f2d240_0 .net "out", 0 0, L_0x5c7c3313f1b0;  alias, 1 drivers
S_0x5c7c32f2cc40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f2ca70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f1b0 .functor NAND 1, L_0x5c7c3313f100, L_0x5c7c3313f100, C4<1>, C4<1>;
v0x5c7c32f2ceb0_0 .net "in_a", 0 0, L_0x5c7c3313f100;  alias, 1 drivers
v0x5c7c32f2cf70_0 .net "in_b", 0 0, L_0x5c7c3313f100;  alias, 1 drivers
v0x5c7c32f2d0c0_0 .net "out", 0 0, L_0x5c7c3313f1b0;  alias, 1 drivers
S_0x5c7c32f2d340 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f28bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f2db10_0 .net "in_a", 0 0, L_0x5c7c3313f420;  alias, 1 drivers
v0x5c7c32f2dbb0_0 .net "out", 0 0, L_0x5c7c3313f4d0;  alias, 1 drivers
S_0x5c7c32f2d5b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f2d340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f4d0 .functor NAND 1, L_0x5c7c3313f420, L_0x5c7c3313f420, C4<1>, C4<1>;
v0x5c7c32f2d820_0 .net "in_a", 0 0, L_0x5c7c3313f420;  alias, 1 drivers
v0x5c7c32f2d8e0_0 .net "in_b", 0 0, L_0x5c7c3313f420;  alias, 1 drivers
v0x5c7c32f2da30_0 .net "out", 0 0, L_0x5c7c3313f4d0;  alias, 1 drivers
S_0x5c7c32f2dcb0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f28bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f2e450_0 .net "in_a", 0 0, L_0x5c7c3313f740;  alias, 1 drivers
v0x5c7c32f2e4f0_0 .net "out", 0 0, L_0x5c7c3313f7f0;  alias, 1 drivers
S_0x5c7c32f2ded0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f2dcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313f7f0 .functor NAND 1, L_0x5c7c3313f740, L_0x5c7c3313f740, C4<1>, C4<1>;
v0x5c7c32f2e140_0 .net "in_a", 0 0, L_0x5c7c3313f740;  alias, 1 drivers
v0x5c7c32f2e200_0 .net "in_b", 0 0, L_0x5c7c3313f740;  alias, 1 drivers
v0x5c7c32f2e350_0 .net "out", 0 0, L_0x5c7c3313f7f0;  alias, 1 drivers
S_0x5c7c32f2f490 .scope module, "mux_gate10" "Mux" 15 17, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f38a10_0 .net "in_a", 0 0, L_0x5c7c33146110;  1 drivers
v0x5c7c32f38ab0_0 .net "in_b", 0 0, L_0x5c7c331483f0;  1 drivers
v0x5c7c32f38bc0_0 .net "out", 0 0, L_0x5c7c33148270;  1 drivers
v0x5c7c32f38c60_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f38d00_0 .net "sel_out", 0 0, L_0x5c7c33146fe0;  1 drivers
v0x5c7c32f38e80_0 .net "temp_a_out", 0 0, L_0x5c7c32f80740;  1 drivers
v0x5c7c32f38f20_0 .net "temp_b_out", 0 0, L_0x5c7c32f808a0;  1 drivers
S_0x5c7c32f2f690 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f2f490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f30700_0 .net "in_a", 0 0, L_0x5c7c33146110;  alias, 1 drivers
v0x5c7c32f307d0_0 .net "in_b", 0 0, L_0x5c7c33146fe0;  alias, 1 drivers
v0x5c7c32f308a0_0 .net "out", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
v0x5c7c32f309c0_0 .net "temp_out", 0 0, L_0x5c7c32f80690;  1 drivers
S_0x5c7c32f2f8e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f2f690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80690 .functor NAND 1, L_0x5c7c33146110, L_0x5c7c33146fe0, C4<1>, C4<1>;
v0x5c7c32f2fb50_0 .net "in_a", 0 0, L_0x5c7c33146110;  alias, 1 drivers
v0x5c7c32f2fc30_0 .net "in_b", 0 0, L_0x5c7c33146fe0;  alias, 1 drivers
v0x5c7c32f2fcf0_0 .net "out", 0 0, L_0x5c7c32f80690;  alias, 1 drivers
S_0x5c7c32f2fe10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f2f690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f30550_0 .net "in_a", 0 0, L_0x5c7c32f80690;  alias, 1 drivers
v0x5c7c32f305f0_0 .net "out", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
S_0x5c7c32f30030 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f2fe10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80740 .functor NAND 1, L_0x5c7c32f80690, L_0x5c7c32f80690, C4<1>, C4<1>;
v0x5c7c32f302a0_0 .net "in_a", 0 0, L_0x5c7c32f80690;  alias, 1 drivers
v0x5c7c32f30360_0 .net "in_b", 0 0, L_0x5c7c32f80690;  alias, 1 drivers
v0x5c7c32f30450_0 .net "out", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
S_0x5c7c32f30a80 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f2f490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f31a90_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f31b30_0 .net "in_b", 0 0, L_0x5c7c331483f0;  alias, 1 drivers
v0x5c7c32f31c20_0 .net "out", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
v0x5c7c32f31d40_0 .net "temp_out", 0 0, L_0x5c7c32f807f0;  1 drivers
S_0x5c7c32f30c60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f30a80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f807f0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c331483f0, C4<1>, C4<1>;
v0x5c7c32f30ed0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f30f90_0 .net "in_b", 0 0, L_0x5c7c331483f0;  alias, 1 drivers
v0x5c7c32f31050_0 .net "out", 0 0, L_0x5c7c32f807f0;  alias, 1 drivers
S_0x5c7c32f31170 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f30a80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f318e0_0 .net "in_a", 0 0, L_0x5c7c32f807f0;  alias, 1 drivers
v0x5c7c32f31980_0 .net "out", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
S_0x5c7c32f31390 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f31170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f808a0 .functor NAND 1, L_0x5c7c32f807f0, L_0x5c7c32f807f0, C4<1>, C4<1>;
v0x5c7c32f31600_0 .net "in_a", 0 0, L_0x5c7c32f807f0;  alias, 1 drivers
v0x5c7c32f316f0_0 .net "in_b", 0 0, L_0x5c7c32f807f0;  alias, 1 drivers
v0x5c7c32f317e0_0 .net "out", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
S_0x5c7c32f31e00 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f2f490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f32500_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f327b0_0 .net "out", 0 0, L_0x5c7c33146fe0;  alias, 1 drivers
S_0x5c7c32f31fd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f31e00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146fe0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f32220_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f322e0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f323a0_0 .net "out", 0 0, L_0x5c7c33146fe0;  alias, 1 drivers
S_0x5c7c32f328b0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f2f490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f38360_0 .net "branch1_out", 0 0, L_0x5c7c32f80ab0;  1 drivers
v0x5c7c32f38490_0 .net "branch2_out", 0 0, L_0x5c7c32f80dd0;  1 drivers
v0x5c7c32f385e0_0 .net "in_a", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
v0x5c7c32f386b0_0 .net "in_b", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
v0x5c7c32f38750_0 .net "out", 0 0, L_0x5c7c33148270;  alias, 1 drivers
v0x5c7c32f387f0_0 .net "temp1_out", 0 0, L_0x5c7c32f80a00;  1 drivers
v0x5c7c32f38890_0 .net "temp2_out", 0 0, L_0x5c7c32f80d20;  1 drivers
v0x5c7c32f38930_0 .net "temp3_out", 0 0, L_0x5c7c33148200;  1 drivers
S_0x5c7c32f32ae0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f328b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f33ba0_0 .net "in_a", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
v0x5c7c32f33c40_0 .net "in_b", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
v0x5c7c32f33d00_0 .net "out", 0 0, L_0x5c7c32f80a00;  alias, 1 drivers
v0x5c7c32f33e20_0 .net "temp_out", 0 0, L_0x5c7c32f80950;  1 drivers
S_0x5c7c32f32d50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f32ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80950 .functor NAND 1, L_0x5c7c32f80740, L_0x5c7c32f80740, C4<1>, C4<1>;
v0x5c7c32f32fc0_0 .net "in_a", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
v0x5c7c32f33080_0 .net "in_b", 0 0, L_0x5c7c32f80740;  alias, 1 drivers
v0x5c7c32f331d0_0 .net "out", 0 0, L_0x5c7c32f80950;  alias, 1 drivers
S_0x5c7c32f332d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f32ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f339f0_0 .net "in_a", 0 0, L_0x5c7c32f80950;  alias, 1 drivers
v0x5c7c32f33a90_0 .net "out", 0 0, L_0x5c7c32f80a00;  alias, 1 drivers
S_0x5c7c32f334a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f332d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80a00 .functor NAND 1, L_0x5c7c32f80950, L_0x5c7c32f80950, C4<1>, C4<1>;
v0x5c7c32f33710_0 .net "in_a", 0 0, L_0x5c7c32f80950;  alias, 1 drivers
v0x5c7c32f33800_0 .net "in_b", 0 0, L_0x5c7c32f80950;  alias, 1 drivers
v0x5c7c32f338f0_0 .net "out", 0 0, L_0x5c7c32f80a00;  alias, 1 drivers
S_0x5c7c32f33f90 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f328b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f34fc0_0 .net "in_a", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
v0x5c7c32f35060_0 .net "in_b", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
v0x5c7c32f35120_0 .net "out", 0 0, L_0x5c7c32f80d20;  alias, 1 drivers
v0x5c7c32f35240_0 .net "temp_out", 0 0, L_0x5c7c32f80c70;  1 drivers
S_0x5c7c32f34170 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f33f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80c70 .functor NAND 1, L_0x5c7c32f808a0, L_0x5c7c32f808a0, C4<1>, C4<1>;
v0x5c7c32f343e0_0 .net "in_a", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
v0x5c7c32f344a0_0 .net "in_b", 0 0, L_0x5c7c32f808a0;  alias, 1 drivers
v0x5c7c32f345f0_0 .net "out", 0 0, L_0x5c7c32f80c70;  alias, 1 drivers
S_0x5c7c32f346f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f33f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f34e10_0 .net "in_a", 0 0, L_0x5c7c32f80c70;  alias, 1 drivers
v0x5c7c32f34eb0_0 .net "out", 0 0, L_0x5c7c32f80d20;  alias, 1 drivers
S_0x5c7c32f348c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f346f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80d20 .functor NAND 1, L_0x5c7c32f80c70, L_0x5c7c32f80c70, C4<1>, C4<1>;
v0x5c7c32f34b30_0 .net "in_a", 0 0, L_0x5c7c32f80c70;  alias, 1 drivers
v0x5c7c32f34c20_0 .net "in_b", 0 0, L_0x5c7c32f80c70;  alias, 1 drivers
v0x5c7c32f34d10_0 .net "out", 0 0, L_0x5c7c32f80d20;  alias, 1 drivers
S_0x5c7c32f353b0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f328b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f363f0_0 .net "in_a", 0 0, L_0x5c7c32f80ab0;  alias, 1 drivers
v0x5c7c32f364c0_0 .net "in_b", 0 0, L_0x5c7c32f80dd0;  alias, 1 drivers
v0x5c7c32f36590_0 .net "out", 0 0, L_0x5c7c33148200;  alias, 1 drivers
v0x5c7c32f366b0_0 .net "temp_out", 0 0, L_0x5c7c33148190;  1 drivers
S_0x5c7c32f35590 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f353b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148190 .functor NAND 1, L_0x5c7c32f80ab0, L_0x5c7c32f80dd0, C4<1>, C4<1>;
v0x5c7c32f357e0_0 .net "in_a", 0 0, L_0x5c7c32f80ab0;  alias, 1 drivers
v0x5c7c32f358c0_0 .net "in_b", 0 0, L_0x5c7c32f80dd0;  alias, 1 drivers
v0x5c7c32f35980_0 .net "out", 0 0, L_0x5c7c33148190;  alias, 1 drivers
S_0x5c7c32f35ad0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f353b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f36240_0 .net "in_a", 0 0, L_0x5c7c33148190;  alias, 1 drivers
v0x5c7c32f362e0_0 .net "out", 0 0, L_0x5c7c33148200;  alias, 1 drivers
S_0x5c7c32f35cf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f35ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148200 .functor NAND 1, L_0x5c7c33148190, L_0x5c7c33148190, C4<1>, C4<1>;
v0x5c7c32f35f60_0 .net "in_a", 0 0, L_0x5c7c33148190;  alias, 1 drivers
v0x5c7c32f36050_0 .net "in_b", 0 0, L_0x5c7c33148190;  alias, 1 drivers
v0x5c7c32f36140_0 .net "out", 0 0, L_0x5c7c33148200;  alias, 1 drivers
S_0x5c7c32f36800 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f328b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f36f30_0 .net "in_a", 0 0, L_0x5c7c32f80a00;  alias, 1 drivers
v0x5c7c32f36fd0_0 .net "out", 0 0, L_0x5c7c32f80ab0;  alias, 1 drivers
S_0x5c7c32f369d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f36800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80ab0 .functor NAND 1, L_0x5c7c32f80a00, L_0x5c7c32f80a00, C4<1>, C4<1>;
v0x5c7c32f36c40_0 .net "in_a", 0 0, L_0x5c7c32f80a00;  alias, 1 drivers
v0x5c7c32f36d00_0 .net "in_b", 0 0, L_0x5c7c32f80a00;  alias, 1 drivers
v0x5c7c32f36e50_0 .net "out", 0 0, L_0x5c7c32f80ab0;  alias, 1 drivers
S_0x5c7c32f370d0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f328b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f378a0_0 .net "in_a", 0 0, L_0x5c7c32f80d20;  alias, 1 drivers
v0x5c7c32f37940_0 .net "out", 0 0, L_0x5c7c32f80dd0;  alias, 1 drivers
S_0x5c7c32f37340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f370d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32f80dd0 .functor NAND 1, L_0x5c7c32f80d20, L_0x5c7c32f80d20, C4<1>, C4<1>;
v0x5c7c32f375b0_0 .net "in_a", 0 0, L_0x5c7c32f80d20;  alias, 1 drivers
v0x5c7c32f37670_0 .net "in_b", 0 0, L_0x5c7c32f80d20;  alias, 1 drivers
v0x5c7c32f377c0_0 .net "out", 0 0, L_0x5c7c32f80dd0;  alias, 1 drivers
S_0x5c7c32f37a40 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f328b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f381e0_0 .net "in_a", 0 0, L_0x5c7c33148200;  alias, 1 drivers
v0x5c7c32f38280_0 .net "out", 0 0, L_0x5c7c33148270;  alias, 1 drivers
S_0x5c7c32f37c60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f37a40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148270 .functor NAND 1, L_0x5c7c33148200, L_0x5c7c33148200, C4<1>, C4<1>;
v0x5c7c32f37ed0_0 .net "in_a", 0 0, L_0x5c7c33148200;  alias, 1 drivers
v0x5c7c32f37f90_0 .net "in_b", 0 0, L_0x5c7c33148200;  alias, 1 drivers
v0x5c7c32f380e0_0 .net "out", 0 0, L_0x5c7c33148270;  alias, 1 drivers
S_0x5c7c32f39110 .scope module, "mux_gate11" "Mux" 15 18, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f42470_0 .net "in_a", 0 0, L_0x5c7c33148ea0;  1 drivers
v0x5c7c32f42510_0 .net "in_b", 0 0, L_0x5c7c33148f40;  1 drivers
v0x5c7c32f42620_0 .net "out", 0 0, L_0x5c7c33148d20;  1 drivers
v0x5c7c32f426c0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f42760_0 .net "sel_out", 0 0, L_0x5c7c33148550;  1 drivers
v0x5c7c32f428e0_0 .net "temp_a_out", 0 0, L_0x5c7c33148630;  1 drivers
v0x5c7c32f42a90_0 .net "temp_b_out", 0 0, L_0x5c7c33148710;  1 drivers
S_0x5c7c32f39310 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f39110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f3a370_0 .net "in_a", 0 0, L_0x5c7c33148ea0;  alias, 1 drivers
v0x5c7c32f3a440_0 .net "in_b", 0 0, L_0x5c7c33148550;  alias, 1 drivers
v0x5c7c32f3a510_0 .net "out", 0 0, L_0x5c7c33148630;  alias, 1 drivers
v0x5c7c32f3a630_0 .net "temp_out", 0 0, L_0x5c7c331485c0;  1 drivers
S_0x5c7c32f39580 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f39310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331485c0 .functor NAND 1, L_0x5c7c33148ea0, L_0x5c7c33148550, C4<1>, C4<1>;
v0x5c7c32f397f0_0 .net "in_a", 0 0, L_0x5c7c33148ea0;  alias, 1 drivers
v0x5c7c32f398d0_0 .net "in_b", 0 0, L_0x5c7c33148550;  alias, 1 drivers
v0x5c7c32f39990_0 .net "out", 0 0, L_0x5c7c331485c0;  alias, 1 drivers
S_0x5c7c32f39ab0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f39310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f3a1f0_0 .net "in_a", 0 0, L_0x5c7c331485c0;  alias, 1 drivers
v0x5c7c32f3a290_0 .net "out", 0 0, L_0x5c7c33148630;  alias, 1 drivers
S_0x5c7c32f39cd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f39ab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148630 .functor NAND 1, L_0x5c7c331485c0, L_0x5c7c331485c0, C4<1>, C4<1>;
v0x5c7c32f39f40_0 .net "in_a", 0 0, L_0x5c7c331485c0;  alias, 1 drivers
v0x5c7c32f3a000_0 .net "in_b", 0 0, L_0x5c7c331485c0;  alias, 1 drivers
v0x5c7c32f3a0f0_0 .net "out", 0 0, L_0x5c7c33148630;  alias, 1 drivers
S_0x5c7c32f3a6f0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f39110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f3b700_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f3b7a0_0 .net "in_b", 0 0, L_0x5c7c33148f40;  alias, 1 drivers
v0x5c7c32f3b890_0 .net "out", 0 0, L_0x5c7c33148710;  alias, 1 drivers
v0x5c7c32f3b9b0_0 .net "temp_out", 0 0, L_0x5c7c331486a0;  1 drivers
S_0x5c7c32f3a8d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f3a6f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331486a0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33148f40, C4<1>, C4<1>;
v0x5c7c32f3ab40_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f3ac00_0 .net "in_b", 0 0, L_0x5c7c33148f40;  alias, 1 drivers
v0x5c7c32f3acc0_0 .net "out", 0 0, L_0x5c7c331486a0;  alias, 1 drivers
S_0x5c7c32f3ade0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f3a6f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f3b550_0 .net "in_a", 0 0, L_0x5c7c331486a0;  alias, 1 drivers
v0x5c7c32f3b5f0_0 .net "out", 0 0, L_0x5c7c33148710;  alias, 1 drivers
S_0x5c7c32f3b000 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f3ade0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148710 .functor NAND 1, L_0x5c7c331486a0, L_0x5c7c331486a0, C4<1>, C4<1>;
v0x5c7c32f3b270_0 .net "in_a", 0 0, L_0x5c7c331486a0;  alias, 1 drivers
v0x5c7c32f3b360_0 .net "in_b", 0 0, L_0x5c7c331486a0;  alias, 1 drivers
v0x5c7c32f3b450_0 .net "out", 0 0, L_0x5c7c33148710;  alias, 1 drivers
S_0x5c7c32f3ba70 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f39110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f3c170_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f3c210_0 .net "out", 0 0, L_0x5c7c33148550;  alias, 1 drivers
S_0x5c7c32f3bc40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f3ba70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148550 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f3be90_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f3bf50_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f3c010_0 .net "out", 0 0, L_0x5c7c33148550;  alias, 1 drivers
S_0x5c7c32f3c310 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f39110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f41dc0_0 .net "branch1_out", 0 0, L_0x5c7c33148860;  1 drivers
v0x5c7c32f41ef0_0 .net "branch2_out", 0 0, L_0x5c7c33148ac0;  1 drivers
v0x5c7c32f42040_0 .net "in_a", 0 0, L_0x5c7c33148630;  alias, 1 drivers
v0x5c7c32f42110_0 .net "in_b", 0 0, L_0x5c7c33148710;  alias, 1 drivers
v0x5c7c32f421b0_0 .net "out", 0 0, L_0x5c7c33148d20;  alias, 1 drivers
v0x5c7c32f42250_0 .net "temp1_out", 0 0, L_0x5c7c331487f0;  1 drivers
v0x5c7c32f422f0_0 .net "temp2_out", 0 0, L_0x5c7c33148a50;  1 drivers
v0x5c7c32f42390_0 .net "temp3_out", 0 0, L_0x5c7c33148cb0;  1 drivers
S_0x5c7c32f3c540 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f3c310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f3d600_0 .net "in_a", 0 0, L_0x5c7c33148630;  alias, 1 drivers
v0x5c7c32f3d6a0_0 .net "in_b", 0 0, L_0x5c7c33148630;  alias, 1 drivers
v0x5c7c32f3d760_0 .net "out", 0 0, L_0x5c7c331487f0;  alias, 1 drivers
v0x5c7c32f3d880_0 .net "temp_out", 0 0, L_0x5c7c33148780;  1 drivers
S_0x5c7c32f3c7b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f3c540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148780 .functor NAND 1, L_0x5c7c33148630, L_0x5c7c33148630, C4<1>, C4<1>;
v0x5c7c32f3ca20_0 .net "in_a", 0 0, L_0x5c7c33148630;  alias, 1 drivers
v0x5c7c32f3cae0_0 .net "in_b", 0 0, L_0x5c7c33148630;  alias, 1 drivers
v0x5c7c32f3cc30_0 .net "out", 0 0, L_0x5c7c33148780;  alias, 1 drivers
S_0x5c7c32f3cd30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f3c540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f3d450_0 .net "in_a", 0 0, L_0x5c7c33148780;  alias, 1 drivers
v0x5c7c32f3d4f0_0 .net "out", 0 0, L_0x5c7c331487f0;  alias, 1 drivers
S_0x5c7c32f3cf00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f3cd30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331487f0 .functor NAND 1, L_0x5c7c33148780, L_0x5c7c33148780, C4<1>, C4<1>;
v0x5c7c32f3d170_0 .net "in_a", 0 0, L_0x5c7c33148780;  alias, 1 drivers
v0x5c7c32f3d260_0 .net "in_b", 0 0, L_0x5c7c33148780;  alias, 1 drivers
v0x5c7c32f3d350_0 .net "out", 0 0, L_0x5c7c331487f0;  alias, 1 drivers
S_0x5c7c32f3d9f0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f3c310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f3ea20_0 .net "in_a", 0 0, L_0x5c7c33148710;  alias, 1 drivers
v0x5c7c32f3eac0_0 .net "in_b", 0 0, L_0x5c7c33148710;  alias, 1 drivers
v0x5c7c32f3eb80_0 .net "out", 0 0, L_0x5c7c33148a50;  alias, 1 drivers
v0x5c7c32f3eca0_0 .net "temp_out", 0 0, L_0x5c7c331489e0;  1 drivers
S_0x5c7c32f3dbd0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f3d9f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331489e0 .functor NAND 1, L_0x5c7c33148710, L_0x5c7c33148710, C4<1>, C4<1>;
v0x5c7c32f3de40_0 .net "in_a", 0 0, L_0x5c7c33148710;  alias, 1 drivers
v0x5c7c32f3df00_0 .net "in_b", 0 0, L_0x5c7c33148710;  alias, 1 drivers
v0x5c7c32f3e050_0 .net "out", 0 0, L_0x5c7c331489e0;  alias, 1 drivers
S_0x5c7c32f3e150 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f3d9f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f3e870_0 .net "in_a", 0 0, L_0x5c7c331489e0;  alias, 1 drivers
v0x5c7c32f3e910_0 .net "out", 0 0, L_0x5c7c33148a50;  alias, 1 drivers
S_0x5c7c32f3e320 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f3e150;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148a50 .functor NAND 1, L_0x5c7c331489e0, L_0x5c7c331489e0, C4<1>, C4<1>;
v0x5c7c32f3e590_0 .net "in_a", 0 0, L_0x5c7c331489e0;  alias, 1 drivers
v0x5c7c32f3e680_0 .net "in_b", 0 0, L_0x5c7c331489e0;  alias, 1 drivers
v0x5c7c32f3e770_0 .net "out", 0 0, L_0x5c7c33148a50;  alias, 1 drivers
S_0x5c7c32f3ee10 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f3c310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f3fe50_0 .net "in_a", 0 0, L_0x5c7c33148860;  alias, 1 drivers
v0x5c7c32f3ff20_0 .net "in_b", 0 0, L_0x5c7c33148ac0;  alias, 1 drivers
v0x5c7c32f3fff0_0 .net "out", 0 0, L_0x5c7c33148cb0;  alias, 1 drivers
v0x5c7c32f40110_0 .net "temp_out", 0 0, L_0x5c7c33148c40;  1 drivers
S_0x5c7c32f3eff0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f3ee10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148c40 .functor NAND 1, L_0x5c7c33148860, L_0x5c7c33148ac0, C4<1>, C4<1>;
v0x5c7c32f3f240_0 .net "in_a", 0 0, L_0x5c7c33148860;  alias, 1 drivers
v0x5c7c32f3f320_0 .net "in_b", 0 0, L_0x5c7c33148ac0;  alias, 1 drivers
v0x5c7c32f3f3e0_0 .net "out", 0 0, L_0x5c7c33148c40;  alias, 1 drivers
S_0x5c7c32f3f530 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f3ee10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f3fca0_0 .net "in_a", 0 0, L_0x5c7c33148c40;  alias, 1 drivers
v0x5c7c32f3fd40_0 .net "out", 0 0, L_0x5c7c33148cb0;  alias, 1 drivers
S_0x5c7c32f3f750 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f3f530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148cb0 .functor NAND 1, L_0x5c7c33148c40, L_0x5c7c33148c40, C4<1>, C4<1>;
v0x5c7c32f3f9c0_0 .net "in_a", 0 0, L_0x5c7c33148c40;  alias, 1 drivers
v0x5c7c32f3fab0_0 .net "in_b", 0 0, L_0x5c7c33148c40;  alias, 1 drivers
v0x5c7c32f3fba0_0 .net "out", 0 0, L_0x5c7c33148cb0;  alias, 1 drivers
S_0x5c7c32f40260 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f3c310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f40990_0 .net "in_a", 0 0, L_0x5c7c331487f0;  alias, 1 drivers
v0x5c7c32f40a30_0 .net "out", 0 0, L_0x5c7c33148860;  alias, 1 drivers
S_0x5c7c32f40430 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f40260;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148860 .functor NAND 1, L_0x5c7c331487f0, L_0x5c7c331487f0, C4<1>, C4<1>;
v0x5c7c32f406a0_0 .net "in_a", 0 0, L_0x5c7c331487f0;  alias, 1 drivers
v0x5c7c32f40760_0 .net "in_b", 0 0, L_0x5c7c331487f0;  alias, 1 drivers
v0x5c7c32f408b0_0 .net "out", 0 0, L_0x5c7c33148860;  alias, 1 drivers
S_0x5c7c32f40b30 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f3c310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f41300_0 .net "in_a", 0 0, L_0x5c7c33148a50;  alias, 1 drivers
v0x5c7c32f413a0_0 .net "out", 0 0, L_0x5c7c33148ac0;  alias, 1 drivers
S_0x5c7c32f40da0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f40b30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148ac0 .functor NAND 1, L_0x5c7c33148a50, L_0x5c7c33148a50, C4<1>, C4<1>;
v0x5c7c32f41010_0 .net "in_a", 0 0, L_0x5c7c33148a50;  alias, 1 drivers
v0x5c7c32f410d0_0 .net "in_b", 0 0, L_0x5c7c33148a50;  alias, 1 drivers
v0x5c7c32f41220_0 .net "out", 0 0, L_0x5c7c33148ac0;  alias, 1 drivers
S_0x5c7c32f414a0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f3c310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f41c40_0 .net "in_a", 0 0, L_0x5c7c33148cb0;  alias, 1 drivers
v0x5c7c32f41ce0_0 .net "out", 0 0, L_0x5c7c33148d20;  alias, 1 drivers
S_0x5c7c32f416c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f414a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33148d20 .functor NAND 1, L_0x5c7c33148cb0, L_0x5c7c33148cb0, C4<1>, C4<1>;
v0x5c7c32f41930_0 .net "in_a", 0 0, L_0x5c7c33148cb0;  alias, 1 drivers
v0x5c7c32f419f0_0 .net "in_b", 0 0, L_0x5c7c33148cb0;  alias, 1 drivers
v0x5c7c32f41b40_0 .net "out", 0 0, L_0x5c7c33148d20;  alias, 1 drivers
S_0x5c7c32f42c80 .scope module, "mux_gate12" "Mux" 15 19, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f4c000_0 .net "in_a", 0 0, L_0x5c7c33149a00;  1 drivers
v0x5c7c32f4c0a0_0 .net "in_b", 0 0, L_0x5c7c33149aa0;  1 drivers
v0x5c7c32f4c1b0_0 .net "out", 0 0, L_0x5c7c33149880;  1 drivers
v0x5c7c32f4c250_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f4c2f0_0 .net "sel_out", 0 0, L_0x5c7c331490b0;  1 drivers
v0x5c7c32f4c470_0 .net "temp_a_out", 0 0, L_0x5c7c33149190;  1 drivers
v0x5c7c32f4c620_0 .net "temp_b_out", 0 0, L_0x5c7c33149270;  1 drivers
S_0x5c7c32f42ed0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f42c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f43f30_0 .net "in_a", 0 0, L_0x5c7c33149a00;  alias, 1 drivers
v0x5c7c32f43fd0_0 .net "in_b", 0 0, L_0x5c7c331490b0;  alias, 1 drivers
v0x5c7c32f440a0_0 .net "out", 0 0, L_0x5c7c33149190;  alias, 1 drivers
v0x5c7c32f441c0_0 .net "temp_out", 0 0, L_0x5c7c33149120;  1 drivers
S_0x5c7c32f43140 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f42ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149120 .functor NAND 1, L_0x5c7c33149a00, L_0x5c7c331490b0, C4<1>, C4<1>;
v0x5c7c32f433b0_0 .net "in_a", 0 0, L_0x5c7c33149a00;  alias, 1 drivers
v0x5c7c32f43490_0 .net "in_b", 0 0, L_0x5c7c331490b0;  alias, 1 drivers
v0x5c7c32f43550_0 .net "out", 0 0, L_0x5c7c33149120;  alias, 1 drivers
S_0x5c7c32f43670 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f42ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f43db0_0 .net "in_a", 0 0, L_0x5c7c33149120;  alias, 1 drivers
v0x5c7c32f43e50_0 .net "out", 0 0, L_0x5c7c33149190;  alias, 1 drivers
S_0x5c7c32f43890 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f43670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149190 .functor NAND 1, L_0x5c7c33149120, L_0x5c7c33149120, C4<1>, C4<1>;
v0x5c7c32f43b00_0 .net "in_a", 0 0, L_0x5c7c33149120;  alias, 1 drivers
v0x5c7c32f43bc0_0 .net "in_b", 0 0, L_0x5c7c33149120;  alias, 1 drivers
v0x5c7c32f43cb0_0 .net "out", 0 0, L_0x5c7c33149190;  alias, 1 drivers
S_0x5c7c32f44280 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f42c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f45290_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f45330_0 .net "in_b", 0 0, L_0x5c7c33149aa0;  alias, 1 drivers
v0x5c7c32f45420_0 .net "out", 0 0, L_0x5c7c33149270;  alias, 1 drivers
v0x5c7c32f45540_0 .net "temp_out", 0 0, L_0x5c7c33149200;  1 drivers
S_0x5c7c32f44460 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f44280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149200 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33149aa0, C4<1>, C4<1>;
v0x5c7c32f446d0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f44790_0 .net "in_b", 0 0, L_0x5c7c33149aa0;  alias, 1 drivers
v0x5c7c32f44850_0 .net "out", 0 0, L_0x5c7c33149200;  alias, 1 drivers
S_0x5c7c32f44970 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f44280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f450e0_0 .net "in_a", 0 0, L_0x5c7c33149200;  alias, 1 drivers
v0x5c7c32f45180_0 .net "out", 0 0, L_0x5c7c33149270;  alias, 1 drivers
S_0x5c7c32f44b90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f44970;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149270 .functor NAND 1, L_0x5c7c33149200, L_0x5c7c33149200, C4<1>, C4<1>;
v0x5c7c32f44e00_0 .net "in_a", 0 0, L_0x5c7c33149200;  alias, 1 drivers
v0x5c7c32f44ef0_0 .net "in_b", 0 0, L_0x5c7c33149200;  alias, 1 drivers
v0x5c7c32f44fe0_0 .net "out", 0 0, L_0x5c7c33149270;  alias, 1 drivers
S_0x5c7c32f45600 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f42c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f45d00_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f45da0_0 .net "out", 0 0, L_0x5c7c331490b0;  alias, 1 drivers
S_0x5c7c32f457d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f45600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331490b0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f45a20_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f45ae0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f45ba0_0 .net "out", 0 0, L_0x5c7c331490b0;  alias, 1 drivers
S_0x5c7c32f45ea0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f42c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f4b950_0 .net "branch1_out", 0 0, L_0x5c7c331493c0;  1 drivers
v0x5c7c32f4ba80_0 .net "branch2_out", 0 0, L_0x5c7c33149620;  1 drivers
v0x5c7c32f4bbd0_0 .net "in_a", 0 0, L_0x5c7c33149190;  alias, 1 drivers
v0x5c7c32f4bca0_0 .net "in_b", 0 0, L_0x5c7c33149270;  alias, 1 drivers
v0x5c7c32f4bd40_0 .net "out", 0 0, L_0x5c7c33149880;  alias, 1 drivers
v0x5c7c32f4bde0_0 .net "temp1_out", 0 0, L_0x5c7c33149350;  1 drivers
v0x5c7c32f4be80_0 .net "temp2_out", 0 0, L_0x5c7c331495b0;  1 drivers
v0x5c7c32f4bf20_0 .net "temp3_out", 0 0, L_0x5c7c33149810;  1 drivers
S_0x5c7c32f460d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f45ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f47190_0 .net "in_a", 0 0, L_0x5c7c33149190;  alias, 1 drivers
v0x5c7c32f47230_0 .net "in_b", 0 0, L_0x5c7c33149190;  alias, 1 drivers
v0x5c7c32f472f0_0 .net "out", 0 0, L_0x5c7c33149350;  alias, 1 drivers
v0x5c7c32f47410_0 .net "temp_out", 0 0, L_0x5c7c331492e0;  1 drivers
S_0x5c7c32f46340 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f460d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331492e0 .functor NAND 1, L_0x5c7c33149190, L_0x5c7c33149190, C4<1>, C4<1>;
v0x5c7c32f465b0_0 .net "in_a", 0 0, L_0x5c7c33149190;  alias, 1 drivers
v0x5c7c32f46670_0 .net "in_b", 0 0, L_0x5c7c33149190;  alias, 1 drivers
v0x5c7c32f467c0_0 .net "out", 0 0, L_0x5c7c331492e0;  alias, 1 drivers
S_0x5c7c32f468c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f460d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f46fe0_0 .net "in_a", 0 0, L_0x5c7c331492e0;  alias, 1 drivers
v0x5c7c32f47080_0 .net "out", 0 0, L_0x5c7c33149350;  alias, 1 drivers
S_0x5c7c32f46a90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f468c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149350 .functor NAND 1, L_0x5c7c331492e0, L_0x5c7c331492e0, C4<1>, C4<1>;
v0x5c7c32f46d00_0 .net "in_a", 0 0, L_0x5c7c331492e0;  alias, 1 drivers
v0x5c7c32f46df0_0 .net "in_b", 0 0, L_0x5c7c331492e0;  alias, 1 drivers
v0x5c7c32f46ee0_0 .net "out", 0 0, L_0x5c7c33149350;  alias, 1 drivers
S_0x5c7c32f47580 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f45ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f485b0_0 .net "in_a", 0 0, L_0x5c7c33149270;  alias, 1 drivers
v0x5c7c32f48650_0 .net "in_b", 0 0, L_0x5c7c33149270;  alias, 1 drivers
v0x5c7c32f48710_0 .net "out", 0 0, L_0x5c7c331495b0;  alias, 1 drivers
v0x5c7c32f48830_0 .net "temp_out", 0 0, L_0x5c7c33149540;  1 drivers
S_0x5c7c32f47760 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f47580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149540 .functor NAND 1, L_0x5c7c33149270, L_0x5c7c33149270, C4<1>, C4<1>;
v0x5c7c32f479d0_0 .net "in_a", 0 0, L_0x5c7c33149270;  alias, 1 drivers
v0x5c7c32f47a90_0 .net "in_b", 0 0, L_0x5c7c33149270;  alias, 1 drivers
v0x5c7c32f47be0_0 .net "out", 0 0, L_0x5c7c33149540;  alias, 1 drivers
S_0x5c7c32f47ce0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f47580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f48400_0 .net "in_a", 0 0, L_0x5c7c33149540;  alias, 1 drivers
v0x5c7c32f484a0_0 .net "out", 0 0, L_0x5c7c331495b0;  alias, 1 drivers
S_0x5c7c32f47eb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f47ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331495b0 .functor NAND 1, L_0x5c7c33149540, L_0x5c7c33149540, C4<1>, C4<1>;
v0x5c7c32f48120_0 .net "in_a", 0 0, L_0x5c7c33149540;  alias, 1 drivers
v0x5c7c32f48210_0 .net "in_b", 0 0, L_0x5c7c33149540;  alias, 1 drivers
v0x5c7c32f48300_0 .net "out", 0 0, L_0x5c7c331495b0;  alias, 1 drivers
S_0x5c7c32f489a0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f45ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f499e0_0 .net "in_a", 0 0, L_0x5c7c331493c0;  alias, 1 drivers
v0x5c7c32f49ab0_0 .net "in_b", 0 0, L_0x5c7c33149620;  alias, 1 drivers
v0x5c7c32f49b80_0 .net "out", 0 0, L_0x5c7c33149810;  alias, 1 drivers
v0x5c7c32f49ca0_0 .net "temp_out", 0 0, L_0x5c7c331497a0;  1 drivers
S_0x5c7c32f48b80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f489a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331497a0 .functor NAND 1, L_0x5c7c331493c0, L_0x5c7c33149620, C4<1>, C4<1>;
v0x5c7c32f48dd0_0 .net "in_a", 0 0, L_0x5c7c331493c0;  alias, 1 drivers
v0x5c7c32f48eb0_0 .net "in_b", 0 0, L_0x5c7c33149620;  alias, 1 drivers
v0x5c7c32f48f70_0 .net "out", 0 0, L_0x5c7c331497a0;  alias, 1 drivers
S_0x5c7c32f490c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f489a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f49830_0 .net "in_a", 0 0, L_0x5c7c331497a0;  alias, 1 drivers
v0x5c7c32f498d0_0 .net "out", 0 0, L_0x5c7c33149810;  alias, 1 drivers
S_0x5c7c32f492e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f490c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149810 .functor NAND 1, L_0x5c7c331497a0, L_0x5c7c331497a0, C4<1>, C4<1>;
v0x5c7c32f49550_0 .net "in_a", 0 0, L_0x5c7c331497a0;  alias, 1 drivers
v0x5c7c32f49640_0 .net "in_b", 0 0, L_0x5c7c331497a0;  alias, 1 drivers
v0x5c7c32f49730_0 .net "out", 0 0, L_0x5c7c33149810;  alias, 1 drivers
S_0x5c7c32f49df0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f45ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f4a520_0 .net "in_a", 0 0, L_0x5c7c33149350;  alias, 1 drivers
v0x5c7c32f4a5c0_0 .net "out", 0 0, L_0x5c7c331493c0;  alias, 1 drivers
S_0x5c7c32f49fc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f49df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331493c0 .functor NAND 1, L_0x5c7c33149350, L_0x5c7c33149350, C4<1>, C4<1>;
v0x5c7c32f4a230_0 .net "in_a", 0 0, L_0x5c7c33149350;  alias, 1 drivers
v0x5c7c32f4a2f0_0 .net "in_b", 0 0, L_0x5c7c33149350;  alias, 1 drivers
v0x5c7c32f4a440_0 .net "out", 0 0, L_0x5c7c331493c0;  alias, 1 drivers
S_0x5c7c32f4a6c0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f45ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f4ae90_0 .net "in_a", 0 0, L_0x5c7c331495b0;  alias, 1 drivers
v0x5c7c32f4af30_0 .net "out", 0 0, L_0x5c7c33149620;  alias, 1 drivers
S_0x5c7c32f4a930 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f4a6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149620 .functor NAND 1, L_0x5c7c331495b0, L_0x5c7c331495b0, C4<1>, C4<1>;
v0x5c7c32f4aba0_0 .net "in_a", 0 0, L_0x5c7c331495b0;  alias, 1 drivers
v0x5c7c32f4ac60_0 .net "in_b", 0 0, L_0x5c7c331495b0;  alias, 1 drivers
v0x5c7c32f4adb0_0 .net "out", 0 0, L_0x5c7c33149620;  alias, 1 drivers
S_0x5c7c32f4b030 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f45ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f4b7d0_0 .net "in_a", 0 0, L_0x5c7c33149810;  alias, 1 drivers
v0x5c7c32f4b870_0 .net "out", 0 0, L_0x5c7c33149880;  alias, 1 drivers
S_0x5c7c32f4b250 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f4b030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149880 .functor NAND 1, L_0x5c7c33149810, L_0x5c7c33149810, C4<1>, C4<1>;
v0x5c7c32f4b4c0_0 .net "in_a", 0 0, L_0x5c7c33149810;  alias, 1 drivers
v0x5c7c32f4b580_0 .net "in_b", 0 0, L_0x5c7c33149810;  alias, 1 drivers
v0x5c7c32f4b6d0_0 .net "out", 0 0, L_0x5c7c33149880;  alias, 1 drivers
S_0x5c7c32f4c810 .scope module, "mux_gate13" "Mux" 15 20, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f55f80_0 .net "in_a", 0 0, L_0x5c7c3314a790;  1 drivers
v0x5c7c32f56020_0 .net "in_b", 0 0, L_0x5c7c3314a830;  1 drivers
v0x5c7c32f56130_0 .net "out", 0 0, L_0x5c7c3314a5d0;  1 drivers
v0x5c7c32f561d0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f56270_0 .net "sel_out", 0 0, L_0x5c7c33149c20;  1 drivers
v0x5c7c32f563f0_0 .net "temp_a_out", 0 0, L_0x5c7c33149d00;  1 drivers
v0x5c7c32f565a0_0 .net "temp_b_out", 0 0, L_0x5c7c33149de0;  1 drivers
S_0x5c7c32f4ca10 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f4c810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f4da70_0 .net "in_a", 0 0, L_0x5c7c3314a790;  alias, 1 drivers
v0x5c7c32f4db40_0 .net "in_b", 0 0, L_0x5c7c33149c20;  alias, 1 drivers
v0x5c7c32f4dc10_0 .net "out", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
v0x5c7c32f4dd30_0 .net "temp_out", 0 0, L_0x5c7c33149c90;  1 drivers
S_0x5c7c32f4cc80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f4ca10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149c90 .functor NAND 1, L_0x5c7c3314a790, L_0x5c7c33149c20, C4<1>, C4<1>;
v0x5c7c32f4cef0_0 .net "in_a", 0 0, L_0x5c7c3314a790;  alias, 1 drivers
v0x5c7c32f4cfd0_0 .net "in_b", 0 0, L_0x5c7c33149c20;  alias, 1 drivers
v0x5c7c32f4d090_0 .net "out", 0 0, L_0x5c7c33149c90;  alias, 1 drivers
S_0x5c7c32f4d1b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f4ca10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f4d8f0_0 .net "in_a", 0 0, L_0x5c7c33149c90;  alias, 1 drivers
v0x5c7c32f4d990_0 .net "out", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
S_0x5c7c32f4d3d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f4d1b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149d00 .functor NAND 1, L_0x5c7c33149c90, L_0x5c7c33149c90, C4<1>, C4<1>;
v0x5c7c32f4d640_0 .net "in_a", 0 0, L_0x5c7c33149c90;  alias, 1 drivers
v0x5c7c32f4d700_0 .net "in_b", 0 0, L_0x5c7c33149c90;  alias, 1 drivers
v0x5c7c32f4d7f0_0 .net "out", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
S_0x5c7c32f4ddf0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f4c810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f4ee00_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f4eea0_0 .net "in_b", 0 0, L_0x5c7c3314a830;  alias, 1 drivers
v0x5c7c32f4ef90_0 .net "out", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
v0x5c7c32f4f0b0_0 .net "temp_out", 0 0, L_0x5c7c33149d70;  1 drivers
S_0x5c7c32f4dfd0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f4ddf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149d70 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314a830, C4<1>, C4<1>;
v0x5c7c32f4e240_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f4e300_0 .net "in_b", 0 0, L_0x5c7c3314a830;  alias, 1 drivers
v0x5c7c32f4e3c0_0 .net "out", 0 0, L_0x5c7c33149d70;  alias, 1 drivers
S_0x5c7c32f4e4e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f4ddf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f4ec50_0 .net "in_a", 0 0, L_0x5c7c33149d70;  alias, 1 drivers
v0x5c7c32f4ecf0_0 .net "out", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
S_0x5c7c32f4e700 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f4e4e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149de0 .functor NAND 1, L_0x5c7c33149d70, L_0x5c7c33149d70, C4<1>, C4<1>;
v0x5c7c32f4e970_0 .net "in_a", 0 0, L_0x5c7c33149d70;  alias, 1 drivers
v0x5c7c32f4ea60_0 .net "in_b", 0 0, L_0x5c7c33149d70;  alias, 1 drivers
v0x5c7c32f4eb50_0 .net "out", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
S_0x5c7c32f4f170 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f4c810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f4fc80_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f4fd20_0 .net "out", 0 0, L_0x5c7c33149c20;  alias, 1 drivers
S_0x5c7c32f4f340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f4f170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149c20 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f4f590_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f4fa60_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f4fb20_0 .net "out", 0 0, L_0x5c7c33149c20;  alias, 1 drivers
S_0x5c7c32f4fe20 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f4c810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f558d0_0 .net "branch1_out", 0 0, L_0x5c7c33149f90;  1 drivers
v0x5c7c32f55a00_0 .net "branch2_out", 0 0, L_0x5c7c3314a2b0;  1 drivers
v0x5c7c32f55b50_0 .net "in_a", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
v0x5c7c32f55c20_0 .net "in_b", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
v0x5c7c32f55cc0_0 .net "out", 0 0, L_0x5c7c3314a5d0;  alias, 1 drivers
v0x5c7c32f55d60_0 .net "temp1_out", 0 0, L_0x5c7c33149ee0;  1 drivers
v0x5c7c32f55e00_0 .net "temp2_out", 0 0, L_0x5c7c3314a200;  1 drivers
v0x5c7c32f55ea0_0 .net "temp3_out", 0 0, L_0x5c7c3314a520;  1 drivers
S_0x5c7c32f50050 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f4fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f51110_0 .net "in_a", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
v0x5c7c32f511b0_0 .net "in_b", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
v0x5c7c32f51270_0 .net "out", 0 0, L_0x5c7c33149ee0;  alias, 1 drivers
v0x5c7c32f51390_0 .net "temp_out", 0 0, L_0x5c7c33149e50;  1 drivers
S_0x5c7c32f502c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f50050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149e50 .functor NAND 1, L_0x5c7c33149d00, L_0x5c7c33149d00, C4<1>, C4<1>;
v0x5c7c32f50530_0 .net "in_a", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
v0x5c7c32f505f0_0 .net "in_b", 0 0, L_0x5c7c33149d00;  alias, 1 drivers
v0x5c7c32f50740_0 .net "out", 0 0, L_0x5c7c33149e50;  alias, 1 drivers
S_0x5c7c32f50840 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f50050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f50f60_0 .net "in_a", 0 0, L_0x5c7c33149e50;  alias, 1 drivers
v0x5c7c32f51000_0 .net "out", 0 0, L_0x5c7c33149ee0;  alias, 1 drivers
S_0x5c7c32f50a10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f50840;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149ee0 .functor NAND 1, L_0x5c7c33149e50, L_0x5c7c33149e50, C4<1>, C4<1>;
v0x5c7c32f50c80_0 .net "in_a", 0 0, L_0x5c7c33149e50;  alias, 1 drivers
v0x5c7c32f50d70_0 .net "in_b", 0 0, L_0x5c7c33149e50;  alias, 1 drivers
v0x5c7c32f50e60_0 .net "out", 0 0, L_0x5c7c33149ee0;  alias, 1 drivers
S_0x5c7c32f51500 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f4fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f52530_0 .net "in_a", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
v0x5c7c32f525d0_0 .net "in_b", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
v0x5c7c32f52690_0 .net "out", 0 0, L_0x5c7c3314a200;  alias, 1 drivers
v0x5c7c32f527b0_0 .net "temp_out", 0 0, L_0x5c7c3314a150;  1 drivers
S_0x5c7c32f516e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f51500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a150 .functor NAND 1, L_0x5c7c33149de0, L_0x5c7c33149de0, C4<1>, C4<1>;
v0x5c7c32f51950_0 .net "in_a", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
v0x5c7c32f51a10_0 .net "in_b", 0 0, L_0x5c7c33149de0;  alias, 1 drivers
v0x5c7c32f51b60_0 .net "out", 0 0, L_0x5c7c3314a150;  alias, 1 drivers
S_0x5c7c32f51c60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f51500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f52380_0 .net "in_a", 0 0, L_0x5c7c3314a150;  alias, 1 drivers
v0x5c7c32f52420_0 .net "out", 0 0, L_0x5c7c3314a200;  alias, 1 drivers
S_0x5c7c32f51e30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f51c60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a200 .functor NAND 1, L_0x5c7c3314a150, L_0x5c7c3314a150, C4<1>, C4<1>;
v0x5c7c32f520a0_0 .net "in_a", 0 0, L_0x5c7c3314a150;  alias, 1 drivers
v0x5c7c32f52190_0 .net "in_b", 0 0, L_0x5c7c3314a150;  alias, 1 drivers
v0x5c7c32f52280_0 .net "out", 0 0, L_0x5c7c3314a200;  alias, 1 drivers
S_0x5c7c32f52920 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f4fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f53960_0 .net "in_a", 0 0, L_0x5c7c33149f90;  alias, 1 drivers
v0x5c7c32f53a30_0 .net "in_b", 0 0, L_0x5c7c3314a2b0;  alias, 1 drivers
v0x5c7c32f53b00_0 .net "out", 0 0, L_0x5c7c3314a520;  alias, 1 drivers
v0x5c7c32f53c20_0 .net "temp_out", 0 0, L_0x5c7c3314a470;  1 drivers
S_0x5c7c32f52b00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f52920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a470 .functor NAND 1, L_0x5c7c33149f90, L_0x5c7c3314a2b0, C4<1>, C4<1>;
v0x5c7c32f52d50_0 .net "in_a", 0 0, L_0x5c7c33149f90;  alias, 1 drivers
v0x5c7c32f52e30_0 .net "in_b", 0 0, L_0x5c7c3314a2b0;  alias, 1 drivers
v0x5c7c32f52ef0_0 .net "out", 0 0, L_0x5c7c3314a470;  alias, 1 drivers
S_0x5c7c32f53040 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f52920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f537b0_0 .net "in_a", 0 0, L_0x5c7c3314a470;  alias, 1 drivers
v0x5c7c32f53850_0 .net "out", 0 0, L_0x5c7c3314a520;  alias, 1 drivers
S_0x5c7c32f53260 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f53040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a520 .functor NAND 1, L_0x5c7c3314a470, L_0x5c7c3314a470, C4<1>, C4<1>;
v0x5c7c32f534d0_0 .net "in_a", 0 0, L_0x5c7c3314a470;  alias, 1 drivers
v0x5c7c32f535c0_0 .net "in_b", 0 0, L_0x5c7c3314a470;  alias, 1 drivers
v0x5c7c32f536b0_0 .net "out", 0 0, L_0x5c7c3314a520;  alias, 1 drivers
S_0x5c7c32f53d70 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f4fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f544a0_0 .net "in_a", 0 0, L_0x5c7c33149ee0;  alias, 1 drivers
v0x5c7c32f54540_0 .net "out", 0 0, L_0x5c7c33149f90;  alias, 1 drivers
S_0x5c7c32f53f40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f53d70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33149f90 .functor NAND 1, L_0x5c7c33149ee0, L_0x5c7c33149ee0, C4<1>, C4<1>;
v0x5c7c32f541b0_0 .net "in_a", 0 0, L_0x5c7c33149ee0;  alias, 1 drivers
v0x5c7c32f54270_0 .net "in_b", 0 0, L_0x5c7c33149ee0;  alias, 1 drivers
v0x5c7c32f543c0_0 .net "out", 0 0, L_0x5c7c33149f90;  alias, 1 drivers
S_0x5c7c32f54640 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f4fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f54e10_0 .net "in_a", 0 0, L_0x5c7c3314a200;  alias, 1 drivers
v0x5c7c32f54eb0_0 .net "out", 0 0, L_0x5c7c3314a2b0;  alias, 1 drivers
S_0x5c7c32f548b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f54640;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a2b0 .functor NAND 1, L_0x5c7c3314a200, L_0x5c7c3314a200, C4<1>, C4<1>;
v0x5c7c32f54b20_0 .net "in_a", 0 0, L_0x5c7c3314a200;  alias, 1 drivers
v0x5c7c32f54be0_0 .net "in_b", 0 0, L_0x5c7c3314a200;  alias, 1 drivers
v0x5c7c32f54d30_0 .net "out", 0 0, L_0x5c7c3314a2b0;  alias, 1 drivers
S_0x5c7c32f54fb0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f4fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f55750_0 .net "in_a", 0 0, L_0x5c7c3314a520;  alias, 1 drivers
v0x5c7c32f557f0_0 .net "out", 0 0, L_0x5c7c3314a5d0;  alias, 1 drivers
S_0x5c7c32f551d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f54fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a5d0 .functor NAND 1, L_0x5c7c3314a520, L_0x5c7c3314a520, C4<1>, C4<1>;
v0x5c7c32f55440_0 .net "in_a", 0 0, L_0x5c7c3314a520;  alias, 1 drivers
v0x5c7c32f55500_0 .net "in_b", 0 0, L_0x5c7c3314a520;  alias, 1 drivers
v0x5c7c32f55650_0 .net "out", 0 0, L_0x5c7c3314a5d0;  alias, 1 drivers
S_0x5c7c32f56790 .scope module, "mux_gate14" "Mux" 15 21, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f5faf0_0 .net "in_a", 0 0, L_0x5c7c3314b690;  1 drivers
v0x5c7c32f5fb90_0 .net "in_b", 0 0, L_0x5c7c3314b730;  1 drivers
v0x5c7c32f5fca0_0 .net "out", 0 0, L_0x5c7c3314b4d0;  1 drivers
v0x5c7c32f5fd40_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f5fde0_0 .net "sel_out", 0 0, L_0x5c7c3314a9c0;  1 drivers
v0x5c7c32f5ff60_0 .net "temp_a_out", 0 0, L_0x5c7c3314ab20;  1 drivers
v0x5c7c32f60110_0 .net "temp_b_out", 0 0, L_0x5c7c3314ac80;  1 drivers
S_0x5c7c32f56990 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f56790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f579f0_0 .net "in_a", 0 0, L_0x5c7c3314b690;  alias, 1 drivers
v0x5c7c32f57ac0_0 .net "in_b", 0 0, L_0x5c7c3314a9c0;  alias, 1 drivers
v0x5c7c32f57b90_0 .net "out", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
v0x5c7c32f57cb0_0 .net "temp_out", 0 0, L_0x5c7c3314aa70;  1 drivers
S_0x5c7c32f56c00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f56990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314aa70 .functor NAND 1, L_0x5c7c3314b690, L_0x5c7c3314a9c0, C4<1>, C4<1>;
v0x5c7c32f56e70_0 .net "in_a", 0 0, L_0x5c7c3314b690;  alias, 1 drivers
v0x5c7c32f56f50_0 .net "in_b", 0 0, L_0x5c7c3314a9c0;  alias, 1 drivers
v0x5c7c32f57010_0 .net "out", 0 0, L_0x5c7c3314aa70;  alias, 1 drivers
S_0x5c7c32f57130 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f56990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f57870_0 .net "in_a", 0 0, L_0x5c7c3314aa70;  alias, 1 drivers
v0x5c7c32f57910_0 .net "out", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
S_0x5c7c32f57350 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f57130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ab20 .functor NAND 1, L_0x5c7c3314aa70, L_0x5c7c3314aa70, C4<1>, C4<1>;
v0x5c7c32f575c0_0 .net "in_a", 0 0, L_0x5c7c3314aa70;  alias, 1 drivers
v0x5c7c32f57680_0 .net "in_b", 0 0, L_0x5c7c3314aa70;  alias, 1 drivers
v0x5c7c32f57770_0 .net "out", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
S_0x5c7c32f57d70 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f56790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f58d80_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f58e20_0 .net "in_b", 0 0, L_0x5c7c3314b730;  alias, 1 drivers
v0x5c7c32f58f10_0 .net "out", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
v0x5c7c32f59030_0 .net "temp_out", 0 0, L_0x5c7c3314abd0;  1 drivers
S_0x5c7c32f57f50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f57d70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314abd0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314b730, C4<1>, C4<1>;
v0x5c7c32f581c0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f58280_0 .net "in_b", 0 0, L_0x5c7c3314b730;  alias, 1 drivers
v0x5c7c32f58340_0 .net "out", 0 0, L_0x5c7c3314abd0;  alias, 1 drivers
S_0x5c7c32f58460 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f57d70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f58bd0_0 .net "in_a", 0 0, L_0x5c7c3314abd0;  alias, 1 drivers
v0x5c7c32f58c70_0 .net "out", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
S_0x5c7c32f58680 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f58460;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ac80 .functor NAND 1, L_0x5c7c3314abd0, L_0x5c7c3314abd0, C4<1>, C4<1>;
v0x5c7c32f588f0_0 .net "in_a", 0 0, L_0x5c7c3314abd0;  alias, 1 drivers
v0x5c7c32f589e0_0 .net "in_b", 0 0, L_0x5c7c3314abd0;  alias, 1 drivers
v0x5c7c32f58ad0_0 .net "out", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
S_0x5c7c32f590f0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f56790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f597f0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f59890_0 .net "out", 0 0, L_0x5c7c3314a9c0;  alias, 1 drivers
S_0x5c7c32f592c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f590f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314a9c0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f59510_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f595d0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f59690_0 .net "out", 0 0, L_0x5c7c3314a9c0;  alias, 1 drivers
S_0x5c7c32f59990 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f56790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f5f440_0 .net "branch1_out", 0 0, L_0x5c7c3314ae90;  1 drivers
v0x5c7c32f5f570_0 .net "branch2_out", 0 0, L_0x5c7c3314b1b0;  1 drivers
v0x5c7c32f5f6c0_0 .net "in_a", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
v0x5c7c32f5f790_0 .net "in_b", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
v0x5c7c32f5f830_0 .net "out", 0 0, L_0x5c7c3314b4d0;  alias, 1 drivers
v0x5c7c32f5f8d0_0 .net "temp1_out", 0 0, L_0x5c7c3314ade0;  1 drivers
v0x5c7c32f5f970_0 .net "temp2_out", 0 0, L_0x5c7c3314b100;  1 drivers
v0x5c7c32f5fa10_0 .net "temp3_out", 0 0, L_0x5c7c3314b420;  1 drivers
S_0x5c7c32f59bc0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f59990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f5ac80_0 .net "in_a", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
v0x5c7c32f5ad20_0 .net "in_b", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
v0x5c7c32f5ade0_0 .net "out", 0 0, L_0x5c7c3314ade0;  alias, 1 drivers
v0x5c7c32f5af00_0 .net "temp_out", 0 0, L_0x5c7c3314ad30;  1 drivers
S_0x5c7c32f59e30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f59bc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ad30 .functor NAND 1, L_0x5c7c3314ab20, L_0x5c7c3314ab20, C4<1>, C4<1>;
v0x5c7c32f5a0a0_0 .net "in_a", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
v0x5c7c32f5a160_0 .net "in_b", 0 0, L_0x5c7c3314ab20;  alias, 1 drivers
v0x5c7c32f5a2b0_0 .net "out", 0 0, L_0x5c7c3314ad30;  alias, 1 drivers
S_0x5c7c32f5a3b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f59bc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f5aad0_0 .net "in_a", 0 0, L_0x5c7c3314ad30;  alias, 1 drivers
v0x5c7c32f5ab70_0 .net "out", 0 0, L_0x5c7c3314ade0;  alias, 1 drivers
S_0x5c7c32f5a580 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f5a3b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ade0 .functor NAND 1, L_0x5c7c3314ad30, L_0x5c7c3314ad30, C4<1>, C4<1>;
v0x5c7c32f5a7f0_0 .net "in_a", 0 0, L_0x5c7c3314ad30;  alias, 1 drivers
v0x5c7c32f5a8e0_0 .net "in_b", 0 0, L_0x5c7c3314ad30;  alias, 1 drivers
v0x5c7c32f5a9d0_0 .net "out", 0 0, L_0x5c7c3314ade0;  alias, 1 drivers
S_0x5c7c32f5b070 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f59990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f5c0a0_0 .net "in_a", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
v0x5c7c32f5c140_0 .net "in_b", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
v0x5c7c32f5c200_0 .net "out", 0 0, L_0x5c7c3314b100;  alias, 1 drivers
v0x5c7c32f5c320_0 .net "temp_out", 0 0, L_0x5c7c3314b050;  1 drivers
S_0x5c7c32f5b250 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f5b070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314b050 .functor NAND 1, L_0x5c7c3314ac80, L_0x5c7c3314ac80, C4<1>, C4<1>;
v0x5c7c32f5b4c0_0 .net "in_a", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
v0x5c7c32f5b580_0 .net "in_b", 0 0, L_0x5c7c3314ac80;  alias, 1 drivers
v0x5c7c32f5b6d0_0 .net "out", 0 0, L_0x5c7c3314b050;  alias, 1 drivers
S_0x5c7c32f5b7d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f5b070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f5bef0_0 .net "in_a", 0 0, L_0x5c7c3314b050;  alias, 1 drivers
v0x5c7c32f5bf90_0 .net "out", 0 0, L_0x5c7c3314b100;  alias, 1 drivers
S_0x5c7c32f5b9a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f5b7d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314b100 .functor NAND 1, L_0x5c7c3314b050, L_0x5c7c3314b050, C4<1>, C4<1>;
v0x5c7c32f5bc10_0 .net "in_a", 0 0, L_0x5c7c3314b050;  alias, 1 drivers
v0x5c7c32f5bd00_0 .net "in_b", 0 0, L_0x5c7c3314b050;  alias, 1 drivers
v0x5c7c32f5bdf0_0 .net "out", 0 0, L_0x5c7c3314b100;  alias, 1 drivers
S_0x5c7c32f5c490 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f59990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f5d4d0_0 .net "in_a", 0 0, L_0x5c7c3314ae90;  alias, 1 drivers
v0x5c7c32f5d5a0_0 .net "in_b", 0 0, L_0x5c7c3314b1b0;  alias, 1 drivers
v0x5c7c32f5d670_0 .net "out", 0 0, L_0x5c7c3314b420;  alias, 1 drivers
v0x5c7c32f5d790_0 .net "temp_out", 0 0, L_0x5c7c3314b370;  1 drivers
S_0x5c7c32f5c670 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f5c490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314b370 .functor NAND 1, L_0x5c7c3314ae90, L_0x5c7c3314b1b0, C4<1>, C4<1>;
v0x5c7c32f5c8c0_0 .net "in_a", 0 0, L_0x5c7c3314ae90;  alias, 1 drivers
v0x5c7c32f5c9a0_0 .net "in_b", 0 0, L_0x5c7c3314b1b0;  alias, 1 drivers
v0x5c7c32f5ca60_0 .net "out", 0 0, L_0x5c7c3314b370;  alias, 1 drivers
S_0x5c7c32f5cbb0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f5c490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f5d320_0 .net "in_a", 0 0, L_0x5c7c3314b370;  alias, 1 drivers
v0x5c7c32f5d3c0_0 .net "out", 0 0, L_0x5c7c3314b420;  alias, 1 drivers
S_0x5c7c32f5cdd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f5cbb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314b420 .functor NAND 1, L_0x5c7c3314b370, L_0x5c7c3314b370, C4<1>, C4<1>;
v0x5c7c32f5d040_0 .net "in_a", 0 0, L_0x5c7c3314b370;  alias, 1 drivers
v0x5c7c32f5d130_0 .net "in_b", 0 0, L_0x5c7c3314b370;  alias, 1 drivers
v0x5c7c32f5d220_0 .net "out", 0 0, L_0x5c7c3314b420;  alias, 1 drivers
S_0x5c7c32f5d8e0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f59990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f5e010_0 .net "in_a", 0 0, L_0x5c7c3314ade0;  alias, 1 drivers
v0x5c7c32f5e0b0_0 .net "out", 0 0, L_0x5c7c3314ae90;  alias, 1 drivers
S_0x5c7c32f5dab0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f5d8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ae90 .functor NAND 1, L_0x5c7c3314ade0, L_0x5c7c3314ade0, C4<1>, C4<1>;
v0x5c7c32f5dd20_0 .net "in_a", 0 0, L_0x5c7c3314ade0;  alias, 1 drivers
v0x5c7c32f5dde0_0 .net "in_b", 0 0, L_0x5c7c3314ade0;  alias, 1 drivers
v0x5c7c32f5df30_0 .net "out", 0 0, L_0x5c7c3314ae90;  alias, 1 drivers
S_0x5c7c32f5e1b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f59990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f5e980_0 .net "in_a", 0 0, L_0x5c7c3314b100;  alias, 1 drivers
v0x5c7c32f5ea20_0 .net "out", 0 0, L_0x5c7c3314b1b0;  alias, 1 drivers
S_0x5c7c32f5e420 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f5e1b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314b1b0 .functor NAND 1, L_0x5c7c3314b100, L_0x5c7c3314b100, C4<1>, C4<1>;
v0x5c7c32f5e690_0 .net "in_a", 0 0, L_0x5c7c3314b100;  alias, 1 drivers
v0x5c7c32f5e750_0 .net "in_b", 0 0, L_0x5c7c3314b100;  alias, 1 drivers
v0x5c7c32f5e8a0_0 .net "out", 0 0, L_0x5c7c3314b1b0;  alias, 1 drivers
S_0x5c7c32f5eb20 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f59990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f5f2c0_0 .net "in_a", 0 0, L_0x5c7c3314b420;  alias, 1 drivers
v0x5c7c32f5f360_0 .net "out", 0 0, L_0x5c7c3314b4d0;  alias, 1 drivers
S_0x5c7c32f5ed40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f5eb20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314b4d0 .functor NAND 1, L_0x5c7c3314b420, L_0x5c7c3314b420, C4<1>, C4<1>;
v0x5c7c32f5efb0_0 .net "in_a", 0 0, L_0x5c7c3314b420;  alias, 1 drivers
v0x5c7c32f5f070_0 .net "in_b", 0 0, L_0x5c7c3314b420;  alias, 1 drivers
v0x5c7c32f5f1c0_0 .net "out", 0 0, L_0x5c7c3314b4d0;  alias, 1 drivers
S_0x5c7c32f60300 .scope module, "mux_gate15" "Mux" 15 22, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f69660_0 .net "in_a", 0 0, L_0x5c7c3314c590;  1 drivers
v0x5c7c32f69700_0 .net "in_b", 0 0, L_0x5c7c3314c630;  1 drivers
v0x5c7c32f69810_0 .net "out", 0 0, L_0x5c7c3314c3d0;  1 drivers
v0x5c7c32f698b0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f69950_0 .net "sel_out", 0 0, L_0x5c7c3314bae0;  1 drivers
v0x5c7c32f69ad0_0 .net "temp_a_out", 0 0, L_0x5c7c3314bc40;  1 drivers
v0x5c7c32f69c80_0 .net "temp_b_out", 0 0, L_0x5c7c3314bda0;  1 drivers
S_0x5c7c32f60500 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f60300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f61560_0 .net "in_a", 0 0, L_0x5c7c3314c590;  alias, 1 drivers
v0x5c7c32f61630_0 .net "in_b", 0 0, L_0x5c7c3314bae0;  alias, 1 drivers
v0x5c7c32f61700_0 .net "out", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
v0x5c7c32f61820_0 .net "temp_out", 0 0, L_0x5c7c3314bb90;  1 drivers
S_0x5c7c32f60770 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f60500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bb90 .functor NAND 1, L_0x5c7c3314c590, L_0x5c7c3314bae0, C4<1>, C4<1>;
v0x5c7c32f609e0_0 .net "in_a", 0 0, L_0x5c7c3314c590;  alias, 1 drivers
v0x5c7c32f60ac0_0 .net "in_b", 0 0, L_0x5c7c3314bae0;  alias, 1 drivers
v0x5c7c32f60b80_0 .net "out", 0 0, L_0x5c7c3314bb90;  alias, 1 drivers
S_0x5c7c32f60ca0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f60500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f613e0_0 .net "in_a", 0 0, L_0x5c7c3314bb90;  alias, 1 drivers
v0x5c7c32f61480_0 .net "out", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
S_0x5c7c32f60ec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f60ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bc40 .functor NAND 1, L_0x5c7c3314bb90, L_0x5c7c3314bb90, C4<1>, C4<1>;
v0x5c7c32f61130_0 .net "in_a", 0 0, L_0x5c7c3314bb90;  alias, 1 drivers
v0x5c7c32f611f0_0 .net "in_b", 0 0, L_0x5c7c3314bb90;  alias, 1 drivers
v0x5c7c32f612e0_0 .net "out", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
S_0x5c7c32f618e0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f60300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f628f0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f62990_0 .net "in_b", 0 0, L_0x5c7c3314c630;  alias, 1 drivers
v0x5c7c32f62a80_0 .net "out", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
v0x5c7c32f62ba0_0 .net "temp_out", 0 0, L_0x5c7c3314bcf0;  1 drivers
S_0x5c7c32f61ac0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f618e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bcf0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c630, C4<1>, C4<1>;
v0x5c7c32f61d30_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f61df0_0 .net "in_b", 0 0, L_0x5c7c3314c630;  alias, 1 drivers
v0x5c7c32f61eb0_0 .net "out", 0 0, L_0x5c7c3314bcf0;  alias, 1 drivers
S_0x5c7c32f61fd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f618e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f62740_0 .net "in_a", 0 0, L_0x5c7c3314bcf0;  alias, 1 drivers
v0x5c7c32f627e0_0 .net "out", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
S_0x5c7c32f621f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f61fd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bda0 .functor NAND 1, L_0x5c7c3314bcf0, L_0x5c7c3314bcf0, C4<1>, C4<1>;
v0x5c7c32f62460_0 .net "in_a", 0 0, L_0x5c7c3314bcf0;  alias, 1 drivers
v0x5c7c32f62550_0 .net "in_b", 0 0, L_0x5c7c3314bcf0;  alias, 1 drivers
v0x5c7c32f62640_0 .net "out", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
S_0x5c7c32f62c60 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f60300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f63360_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f63400_0 .net "out", 0 0, L_0x5c7c3314bae0;  alias, 1 drivers
S_0x5c7c32f62e30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f62c60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bae0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f63080_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f63140_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f63200_0 .net "out", 0 0, L_0x5c7c3314bae0;  alias, 1 drivers
S_0x5c7c32f63500 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f60300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f68fb0_0 .net "branch1_out", 0 0, L_0x5c7c3314bfb0;  1 drivers
v0x5c7c32f690e0_0 .net "branch2_out", 0 0, L_0x5c7c3314c1c0;  1 drivers
v0x5c7c32f69230_0 .net "in_a", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
v0x5c7c32f69300_0 .net "in_b", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
v0x5c7c32f693a0_0 .net "out", 0 0, L_0x5c7c3314c3d0;  alias, 1 drivers
v0x5c7c32f69440_0 .net "temp1_out", 0 0, L_0x5c7c3314bf00;  1 drivers
v0x5c7c32f694e0_0 .net "temp2_out", 0 0, L_0x5c7c3314c110;  1 drivers
v0x5c7c32f69580_0 .net "temp3_out", 0 0, L_0x5c7c3314c320;  1 drivers
S_0x5c7c32f63730 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f63500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f647f0_0 .net "in_a", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
v0x5c7c32f64890_0 .net "in_b", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
v0x5c7c32f64950_0 .net "out", 0 0, L_0x5c7c3314bf00;  alias, 1 drivers
v0x5c7c32f64a70_0 .net "temp_out", 0 0, L_0x5c7c3314be50;  1 drivers
S_0x5c7c32f639a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f63730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314be50 .functor NAND 1, L_0x5c7c3314bc40, L_0x5c7c3314bc40, C4<1>, C4<1>;
v0x5c7c32f63c10_0 .net "in_a", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
v0x5c7c32f63cd0_0 .net "in_b", 0 0, L_0x5c7c3314bc40;  alias, 1 drivers
v0x5c7c32f63e20_0 .net "out", 0 0, L_0x5c7c3314be50;  alias, 1 drivers
S_0x5c7c32f63f20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f63730;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f64640_0 .net "in_a", 0 0, L_0x5c7c3314be50;  alias, 1 drivers
v0x5c7c32f646e0_0 .net "out", 0 0, L_0x5c7c3314bf00;  alias, 1 drivers
S_0x5c7c32f640f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f63f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bf00 .functor NAND 1, L_0x5c7c3314be50, L_0x5c7c3314be50, C4<1>, C4<1>;
v0x5c7c32f64360_0 .net "in_a", 0 0, L_0x5c7c3314be50;  alias, 1 drivers
v0x5c7c32f64450_0 .net "in_b", 0 0, L_0x5c7c3314be50;  alias, 1 drivers
v0x5c7c32f64540_0 .net "out", 0 0, L_0x5c7c3314bf00;  alias, 1 drivers
S_0x5c7c32f64be0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f63500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f65c10_0 .net "in_a", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
v0x5c7c32f65cb0_0 .net "in_b", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
v0x5c7c32f65d70_0 .net "out", 0 0, L_0x5c7c3314c110;  alias, 1 drivers
v0x5c7c32f65e90_0 .net "temp_out", 0 0, L_0x5c7c3314c060;  1 drivers
S_0x5c7c32f64dc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f64be0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c060 .functor NAND 1, L_0x5c7c3314bda0, L_0x5c7c3314bda0, C4<1>, C4<1>;
v0x5c7c32f65030_0 .net "in_a", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
v0x5c7c32f650f0_0 .net "in_b", 0 0, L_0x5c7c3314bda0;  alias, 1 drivers
v0x5c7c32f65240_0 .net "out", 0 0, L_0x5c7c3314c060;  alias, 1 drivers
S_0x5c7c32f65340 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f64be0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f65a60_0 .net "in_a", 0 0, L_0x5c7c3314c060;  alias, 1 drivers
v0x5c7c32f65b00_0 .net "out", 0 0, L_0x5c7c3314c110;  alias, 1 drivers
S_0x5c7c32f65510 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f65340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c110 .functor NAND 1, L_0x5c7c3314c060, L_0x5c7c3314c060, C4<1>, C4<1>;
v0x5c7c32f65780_0 .net "in_a", 0 0, L_0x5c7c3314c060;  alias, 1 drivers
v0x5c7c32f65870_0 .net "in_b", 0 0, L_0x5c7c3314c060;  alias, 1 drivers
v0x5c7c32f65960_0 .net "out", 0 0, L_0x5c7c3314c110;  alias, 1 drivers
S_0x5c7c32f66000 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f63500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f67040_0 .net "in_a", 0 0, L_0x5c7c3314bfb0;  alias, 1 drivers
v0x5c7c32f67110_0 .net "in_b", 0 0, L_0x5c7c3314c1c0;  alias, 1 drivers
v0x5c7c32f671e0_0 .net "out", 0 0, L_0x5c7c3314c320;  alias, 1 drivers
v0x5c7c32f67300_0 .net "temp_out", 0 0, L_0x5c7c3314c270;  1 drivers
S_0x5c7c32f661e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f66000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c270 .functor NAND 1, L_0x5c7c3314bfb0, L_0x5c7c3314c1c0, C4<1>, C4<1>;
v0x5c7c32f66430_0 .net "in_a", 0 0, L_0x5c7c3314bfb0;  alias, 1 drivers
v0x5c7c32f66510_0 .net "in_b", 0 0, L_0x5c7c3314c1c0;  alias, 1 drivers
v0x5c7c32f665d0_0 .net "out", 0 0, L_0x5c7c3314c270;  alias, 1 drivers
S_0x5c7c32f66720 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f66000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f66e90_0 .net "in_a", 0 0, L_0x5c7c3314c270;  alias, 1 drivers
v0x5c7c32f66f30_0 .net "out", 0 0, L_0x5c7c3314c320;  alias, 1 drivers
S_0x5c7c32f66940 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f66720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c320 .functor NAND 1, L_0x5c7c3314c270, L_0x5c7c3314c270, C4<1>, C4<1>;
v0x5c7c32f66bb0_0 .net "in_a", 0 0, L_0x5c7c3314c270;  alias, 1 drivers
v0x5c7c32f66ca0_0 .net "in_b", 0 0, L_0x5c7c3314c270;  alias, 1 drivers
v0x5c7c32f66d90_0 .net "out", 0 0, L_0x5c7c3314c320;  alias, 1 drivers
S_0x5c7c32f67450 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f63500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f67b80_0 .net "in_a", 0 0, L_0x5c7c3314bf00;  alias, 1 drivers
v0x5c7c32f67c20_0 .net "out", 0 0, L_0x5c7c3314bfb0;  alias, 1 drivers
S_0x5c7c32f67620 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f67450;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314bfb0 .functor NAND 1, L_0x5c7c3314bf00, L_0x5c7c3314bf00, C4<1>, C4<1>;
v0x5c7c32f67890_0 .net "in_a", 0 0, L_0x5c7c3314bf00;  alias, 1 drivers
v0x5c7c32f67950_0 .net "in_b", 0 0, L_0x5c7c3314bf00;  alias, 1 drivers
v0x5c7c32f67aa0_0 .net "out", 0 0, L_0x5c7c3314bfb0;  alias, 1 drivers
S_0x5c7c32f67d20 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f63500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f684f0_0 .net "in_a", 0 0, L_0x5c7c3314c110;  alias, 1 drivers
v0x5c7c32f68590_0 .net "out", 0 0, L_0x5c7c3314c1c0;  alias, 1 drivers
S_0x5c7c32f67f90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f67d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c1c0 .functor NAND 1, L_0x5c7c3314c110, L_0x5c7c3314c110, C4<1>, C4<1>;
v0x5c7c32f68200_0 .net "in_a", 0 0, L_0x5c7c3314c110;  alias, 1 drivers
v0x5c7c32f682c0_0 .net "in_b", 0 0, L_0x5c7c3314c110;  alias, 1 drivers
v0x5c7c32f68410_0 .net "out", 0 0, L_0x5c7c3314c1c0;  alias, 1 drivers
S_0x5c7c32f68690 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f63500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f68e30_0 .net "in_a", 0 0, L_0x5c7c3314c320;  alias, 1 drivers
v0x5c7c32f68ed0_0 .net "out", 0 0, L_0x5c7c3314c3d0;  alias, 1 drivers
S_0x5c7c32f688b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f68690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c3d0 .functor NAND 1, L_0x5c7c3314c320, L_0x5c7c3314c320, C4<1>, C4<1>;
v0x5c7c32f68b20_0 .net "in_a", 0 0, L_0x5c7c3314c320;  alias, 1 drivers
v0x5c7c32f68be0_0 .net "in_b", 0 0, L_0x5c7c3314c320;  alias, 1 drivers
v0x5c7c32f68d30_0 .net "out", 0 0, L_0x5c7c3314c3d0;  alias, 1 drivers
S_0x5c7c32f69e70 .scope module, "mux_gate2" "Mux" 15 9, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f73210_0 .net "in_a", 0 0, L_0x5c7c331407a0;  1 drivers
v0x5c7c32f732b0_0 .net "in_b", 0 0, L_0x5c7c33140840;  1 drivers
v0x5c7c32f733c0_0 .net "out", 0 0, L_0x5c7c331405e0;  1 drivers
v0x5c7c32f73460_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f73500_0 .net "sel_out", 0 0, L_0x5c7c3313faf0;  1 drivers
v0x5c7c32f73680_0 .net "temp_a_out", 0 0, L_0x5c7c3313fc30;  1 drivers
v0x5c7c32f73830_0 .net "temp_b_out", 0 0, L_0x5c7c3313fd90;  1 drivers
S_0x5c7c32f6a070 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f69e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f6b080_0 .net "in_a", 0 0, L_0x5c7c331407a0;  alias, 1 drivers
v0x5c7c32f6b150_0 .net "in_b", 0 0, L_0x5c7c3313faf0;  alias, 1 drivers
v0x5c7c32f6b220_0 .net "out", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
v0x5c7c32f6b340_0 .net "temp_out", 0 0, L_0x5c7c3313fb80;  1 drivers
S_0x5c7c32f6a290 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f6a070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313fb80 .functor NAND 1, L_0x5c7c331407a0, L_0x5c7c3313faf0, C4<1>, C4<1>;
v0x5c7c32f6a500_0 .net "in_a", 0 0, L_0x5c7c331407a0;  alias, 1 drivers
v0x5c7c32f6a5e0_0 .net "in_b", 0 0, L_0x5c7c3313faf0;  alias, 1 drivers
v0x5c7c32f6a6a0_0 .net "out", 0 0, L_0x5c7c3313fb80;  alias, 1 drivers
S_0x5c7c32f6a7c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f6a070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f6af00_0 .net "in_a", 0 0, L_0x5c7c3313fb80;  alias, 1 drivers
v0x5c7c32f6afa0_0 .net "out", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
S_0x5c7c32f6a9e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f6a7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313fc30 .functor NAND 1, L_0x5c7c3313fb80, L_0x5c7c3313fb80, C4<1>, C4<1>;
v0x5c7c32f6ac50_0 .net "in_a", 0 0, L_0x5c7c3313fb80;  alias, 1 drivers
v0x5c7c32f6ad10_0 .net "in_b", 0 0, L_0x5c7c3313fb80;  alias, 1 drivers
v0x5c7c32f6ae00_0 .net "out", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
S_0x5c7c32f6b400 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f69e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f6c410_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f6c4b0_0 .net "in_b", 0 0, L_0x5c7c33140840;  alias, 1 drivers
v0x5c7c32f6c5a0_0 .net "out", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
v0x5c7c32f6c6c0_0 .net "temp_out", 0 0, L_0x5c7c3313fce0;  1 drivers
S_0x5c7c32f6b5e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f6b400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313fce0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33140840, C4<1>, C4<1>;
v0x5c7c32f6b850_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f6b910_0 .net "in_b", 0 0, L_0x5c7c33140840;  alias, 1 drivers
v0x5c7c32f6b9d0_0 .net "out", 0 0, L_0x5c7c3313fce0;  alias, 1 drivers
S_0x5c7c32f6baf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f6b400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f6c260_0 .net "in_a", 0 0, L_0x5c7c3313fce0;  alias, 1 drivers
v0x5c7c32f6c300_0 .net "out", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
S_0x5c7c32f6bd10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f6baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313fd90 .functor NAND 1, L_0x5c7c3313fce0, L_0x5c7c3313fce0, C4<1>, C4<1>;
v0x5c7c32f6bf80_0 .net "in_a", 0 0, L_0x5c7c3313fce0;  alias, 1 drivers
v0x5c7c32f6c070_0 .net "in_b", 0 0, L_0x5c7c3313fce0;  alias, 1 drivers
v0x5c7c32f6c160_0 .net "out", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
S_0x5c7c32f6c810 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f69e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f6cf10_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f6cfb0_0 .net "out", 0 0, L_0x5c7c3313faf0;  alias, 1 drivers
S_0x5c7c32f6c9e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f6c810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313faf0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f6cc30_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f6ccf0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f6cdb0_0 .net "out", 0 0, L_0x5c7c3313faf0;  alias, 1 drivers
S_0x5c7c32f6d0b0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f69e70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f72b60_0 .net "branch1_out", 0 0, L_0x5c7c3313ffa0;  1 drivers
v0x5c7c32f72c90_0 .net "branch2_out", 0 0, L_0x5c7c331402c0;  1 drivers
v0x5c7c32f72de0_0 .net "in_a", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
v0x5c7c32f72eb0_0 .net "in_b", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
v0x5c7c32f72f50_0 .net "out", 0 0, L_0x5c7c331405e0;  alias, 1 drivers
v0x5c7c32f72ff0_0 .net "temp1_out", 0 0, L_0x5c7c3313fef0;  1 drivers
v0x5c7c32f73090_0 .net "temp2_out", 0 0, L_0x5c7c33140210;  1 drivers
v0x5c7c32f73130_0 .net "temp3_out", 0 0, L_0x5c7c33140530;  1 drivers
S_0x5c7c32f6d2e0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f6d0b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f6e3a0_0 .net "in_a", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
v0x5c7c32f6e440_0 .net "in_b", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
v0x5c7c32f6e500_0 .net "out", 0 0, L_0x5c7c3313fef0;  alias, 1 drivers
v0x5c7c32f6e620_0 .net "temp_out", 0 0, L_0x5c7c3313fe40;  1 drivers
S_0x5c7c32f6d550 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f6d2e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313fe40 .functor NAND 1, L_0x5c7c3313fc30, L_0x5c7c3313fc30, C4<1>, C4<1>;
v0x5c7c32f6d7c0_0 .net "in_a", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
v0x5c7c32f6d880_0 .net "in_b", 0 0, L_0x5c7c3313fc30;  alias, 1 drivers
v0x5c7c32f6d9d0_0 .net "out", 0 0, L_0x5c7c3313fe40;  alias, 1 drivers
S_0x5c7c32f6dad0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f6d2e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f6e1f0_0 .net "in_a", 0 0, L_0x5c7c3313fe40;  alias, 1 drivers
v0x5c7c32f6e290_0 .net "out", 0 0, L_0x5c7c3313fef0;  alias, 1 drivers
S_0x5c7c32f6dca0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f6dad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313fef0 .functor NAND 1, L_0x5c7c3313fe40, L_0x5c7c3313fe40, C4<1>, C4<1>;
v0x5c7c32f6df10_0 .net "in_a", 0 0, L_0x5c7c3313fe40;  alias, 1 drivers
v0x5c7c32f6e000_0 .net "in_b", 0 0, L_0x5c7c3313fe40;  alias, 1 drivers
v0x5c7c32f6e0f0_0 .net "out", 0 0, L_0x5c7c3313fef0;  alias, 1 drivers
S_0x5c7c32f6e790 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f6d0b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f6f7c0_0 .net "in_a", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
v0x5c7c32f6f860_0 .net "in_b", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
v0x5c7c32f6f920_0 .net "out", 0 0, L_0x5c7c33140210;  alias, 1 drivers
v0x5c7c32f6fa40_0 .net "temp_out", 0 0, L_0x5c7c33140160;  1 drivers
S_0x5c7c32f6e970 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f6e790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140160 .functor NAND 1, L_0x5c7c3313fd90, L_0x5c7c3313fd90, C4<1>, C4<1>;
v0x5c7c32f6ebe0_0 .net "in_a", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
v0x5c7c32f6eca0_0 .net "in_b", 0 0, L_0x5c7c3313fd90;  alias, 1 drivers
v0x5c7c32f6edf0_0 .net "out", 0 0, L_0x5c7c33140160;  alias, 1 drivers
S_0x5c7c32f6eef0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f6e790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f6f610_0 .net "in_a", 0 0, L_0x5c7c33140160;  alias, 1 drivers
v0x5c7c32f6f6b0_0 .net "out", 0 0, L_0x5c7c33140210;  alias, 1 drivers
S_0x5c7c32f6f0c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f6eef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140210 .functor NAND 1, L_0x5c7c33140160, L_0x5c7c33140160, C4<1>, C4<1>;
v0x5c7c32f6f330_0 .net "in_a", 0 0, L_0x5c7c33140160;  alias, 1 drivers
v0x5c7c32f6f420_0 .net "in_b", 0 0, L_0x5c7c33140160;  alias, 1 drivers
v0x5c7c32f6f510_0 .net "out", 0 0, L_0x5c7c33140210;  alias, 1 drivers
S_0x5c7c32f6fbb0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f6d0b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f70bf0_0 .net "in_a", 0 0, L_0x5c7c3313ffa0;  alias, 1 drivers
v0x5c7c32f70cc0_0 .net "in_b", 0 0, L_0x5c7c331402c0;  alias, 1 drivers
v0x5c7c32f70d90_0 .net "out", 0 0, L_0x5c7c33140530;  alias, 1 drivers
v0x5c7c32f70eb0_0 .net "temp_out", 0 0, L_0x5c7c33140480;  1 drivers
S_0x5c7c32f6fd90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f6fbb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140480 .functor NAND 1, L_0x5c7c3313ffa0, L_0x5c7c331402c0, C4<1>, C4<1>;
v0x5c7c32f6ffe0_0 .net "in_a", 0 0, L_0x5c7c3313ffa0;  alias, 1 drivers
v0x5c7c32f700c0_0 .net "in_b", 0 0, L_0x5c7c331402c0;  alias, 1 drivers
v0x5c7c32f70180_0 .net "out", 0 0, L_0x5c7c33140480;  alias, 1 drivers
S_0x5c7c32f702d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f6fbb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f70a40_0 .net "in_a", 0 0, L_0x5c7c33140480;  alias, 1 drivers
v0x5c7c32f70ae0_0 .net "out", 0 0, L_0x5c7c33140530;  alias, 1 drivers
S_0x5c7c32f704f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f702d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140530 .functor NAND 1, L_0x5c7c33140480, L_0x5c7c33140480, C4<1>, C4<1>;
v0x5c7c32f70760_0 .net "in_a", 0 0, L_0x5c7c33140480;  alias, 1 drivers
v0x5c7c32f70850_0 .net "in_b", 0 0, L_0x5c7c33140480;  alias, 1 drivers
v0x5c7c32f70940_0 .net "out", 0 0, L_0x5c7c33140530;  alias, 1 drivers
S_0x5c7c32f71000 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f6d0b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f71730_0 .net "in_a", 0 0, L_0x5c7c3313fef0;  alias, 1 drivers
v0x5c7c32f717d0_0 .net "out", 0 0, L_0x5c7c3313ffa0;  alias, 1 drivers
S_0x5c7c32f711d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f71000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3313ffa0 .functor NAND 1, L_0x5c7c3313fef0, L_0x5c7c3313fef0, C4<1>, C4<1>;
v0x5c7c32f71440_0 .net "in_a", 0 0, L_0x5c7c3313fef0;  alias, 1 drivers
v0x5c7c32f71500_0 .net "in_b", 0 0, L_0x5c7c3313fef0;  alias, 1 drivers
v0x5c7c32f71650_0 .net "out", 0 0, L_0x5c7c3313ffa0;  alias, 1 drivers
S_0x5c7c32f718d0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f6d0b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f720a0_0 .net "in_a", 0 0, L_0x5c7c33140210;  alias, 1 drivers
v0x5c7c32f72140_0 .net "out", 0 0, L_0x5c7c331402c0;  alias, 1 drivers
S_0x5c7c32f71b40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f718d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331402c0 .functor NAND 1, L_0x5c7c33140210, L_0x5c7c33140210, C4<1>, C4<1>;
v0x5c7c32f71db0_0 .net "in_a", 0 0, L_0x5c7c33140210;  alias, 1 drivers
v0x5c7c32f71e70_0 .net "in_b", 0 0, L_0x5c7c33140210;  alias, 1 drivers
v0x5c7c32f71fc0_0 .net "out", 0 0, L_0x5c7c331402c0;  alias, 1 drivers
S_0x5c7c32f72240 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f6d0b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f729e0_0 .net "in_a", 0 0, L_0x5c7c33140530;  alias, 1 drivers
v0x5c7c32f72a80_0 .net "out", 0 0, L_0x5c7c331405e0;  alias, 1 drivers
S_0x5c7c32f72460 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f72240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331405e0 .functor NAND 1, L_0x5c7c33140530, L_0x5c7c33140530, C4<1>, C4<1>;
v0x5c7c32f726d0_0 .net "in_a", 0 0, L_0x5c7c33140530;  alias, 1 drivers
v0x5c7c32f72790_0 .net "in_b", 0 0, L_0x5c7c33140530;  alias, 1 drivers
v0x5c7c32f728e0_0 .net "out", 0 0, L_0x5c7c331405e0;  alias, 1 drivers
S_0x5c7c32f73a20 .scope module, "mux_gate3" "Mux" 15 10, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f7cd80_0 .net "in_a", 0 0, L_0x5c7c331415f0;  1 drivers
v0x5c7c32f7ce20_0 .net "in_b", 0 0, L_0x5c7c33141690;  1 drivers
v0x5c7c32f7cf30_0 .net "out", 0 0, L_0x5c7c33141430;  1 drivers
v0x5c7c32f7cfd0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f7d070_0 .net "sel_out", 0 0, L_0x5c7c33140920;  1 drivers
v0x5c7c32f7d1f0_0 .net "temp_a_out", 0 0, L_0x5c7c33140a80;  1 drivers
v0x5c7c32f7d3a0_0 .net "temp_b_out", 0 0, L_0x5c7c33140be0;  1 drivers
S_0x5c7c32f73c20 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f73a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f74c80_0 .net "in_a", 0 0, L_0x5c7c331415f0;  alias, 1 drivers
v0x5c7c32f74d50_0 .net "in_b", 0 0, L_0x5c7c33140920;  alias, 1 drivers
v0x5c7c32f74e20_0 .net "out", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
v0x5c7c32f74f40_0 .net "temp_out", 0 0, L_0x5c7c331409d0;  1 drivers
S_0x5c7c32f73e90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f73c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331409d0 .functor NAND 1, L_0x5c7c331415f0, L_0x5c7c33140920, C4<1>, C4<1>;
v0x5c7c32f74100_0 .net "in_a", 0 0, L_0x5c7c331415f0;  alias, 1 drivers
v0x5c7c32f741e0_0 .net "in_b", 0 0, L_0x5c7c33140920;  alias, 1 drivers
v0x5c7c32f742a0_0 .net "out", 0 0, L_0x5c7c331409d0;  alias, 1 drivers
S_0x5c7c32f743c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f73c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f74b00_0 .net "in_a", 0 0, L_0x5c7c331409d0;  alias, 1 drivers
v0x5c7c32f74ba0_0 .net "out", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
S_0x5c7c32f745e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f743c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140a80 .functor NAND 1, L_0x5c7c331409d0, L_0x5c7c331409d0, C4<1>, C4<1>;
v0x5c7c32f74850_0 .net "in_a", 0 0, L_0x5c7c331409d0;  alias, 1 drivers
v0x5c7c32f74910_0 .net "in_b", 0 0, L_0x5c7c331409d0;  alias, 1 drivers
v0x5c7c32f74a00_0 .net "out", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
S_0x5c7c32f75000 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f73a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f76010_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f760b0_0 .net "in_b", 0 0, L_0x5c7c33141690;  alias, 1 drivers
v0x5c7c32f761a0_0 .net "out", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
v0x5c7c32f762c0_0 .net "temp_out", 0 0, L_0x5c7c33140b30;  1 drivers
S_0x5c7c32f751e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f75000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140b30 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33141690, C4<1>, C4<1>;
v0x5c7c32f75450_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f75510_0 .net "in_b", 0 0, L_0x5c7c33141690;  alias, 1 drivers
v0x5c7c32f755d0_0 .net "out", 0 0, L_0x5c7c33140b30;  alias, 1 drivers
S_0x5c7c32f756f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f75000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f75e60_0 .net "in_a", 0 0, L_0x5c7c33140b30;  alias, 1 drivers
v0x5c7c32f75f00_0 .net "out", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
S_0x5c7c32f75910 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f756f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140be0 .functor NAND 1, L_0x5c7c33140b30, L_0x5c7c33140b30, C4<1>, C4<1>;
v0x5c7c32f75b80_0 .net "in_a", 0 0, L_0x5c7c33140b30;  alias, 1 drivers
v0x5c7c32f75c70_0 .net "in_b", 0 0, L_0x5c7c33140b30;  alias, 1 drivers
v0x5c7c32f75d60_0 .net "out", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
S_0x5c7c32f76380 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f73a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f76a80_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f76b20_0 .net "out", 0 0, L_0x5c7c33140920;  alias, 1 drivers
S_0x5c7c32f76550 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f76380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140920 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f767a0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f76860_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f76920_0 .net "out", 0 0, L_0x5c7c33140920;  alias, 1 drivers
S_0x5c7c32f76c20 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f73a20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f7c6d0_0 .net "branch1_out", 0 0, L_0x5c7c33140df0;  1 drivers
v0x5c7c32f7c800_0 .net "branch2_out", 0 0, L_0x5c7c33141110;  1 drivers
v0x5c7c32f7c950_0 .net "in_a", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
v0x5c7c32f7ca20_0 .net "in_b", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
v0x5c7c32f7cac0_0 .net "out", 0 0, L_0x5c7c33141430;  alias, 1 drivers
v0x5c7c32f7cb60_0 .net "temp1_out", 0 0, L_0x5c7c33140d40;  1 drivers
v0x5c7c32f7cc00_0 .net "temp2_out", 0 0, L_0x5c7c33141060;  1 drivers
v0x5c7c32f7cca0_0 .net "temp3_out", 0 0, L_0x5c7c33141380;  1 drivers
S_0x5c7c32f76e50 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f76c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f77f10_0 .net "in_a", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
v0x5c7c32f77fb0_0 .net "in_b", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
v0x5c7c32f78070_0 .net "out", 0 0, L_0x5c7c33140d40;  alias, 1 drivers
v0x5c7c32f78190_0 .net "temp_out", 0 0, L_0x5c7c33140c90;  1 drivers
S_0x5c7c32f770c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f76e50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140c90 .functor NAND 1, L_0x5c7c33140a80, L_0x5c7c33140a80, C4<1>, C4<1>;
v0x5c7c32f77330_0 .net "in_a", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
v0x5c7c32f773f0_0 .net "in_b", 0 0, L_0x5c7c33140a80;  alias, 1 drivers
v0x5c7c32f77540_0 .net "out", 0 0, L_0x5c7c33140c90;  alias, 1 drivers
S_0x5c7c32f77640 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f76e50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f77d60_0 .net "in_a", 0 0, L_0x5c7c33140c90;  alias, 1 drivers
v0x5c7c32f77e00_0 .net "out", 0 0, L_0x5c7c33140d40;  alias, 1 drivers
S_0x5c7c32f77810 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f77640;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140d40 .functor NAND 1, L_0x5c7c33140c90, L_0x5c7c33140c90, C4<1>, C4<1>;
v0x5c7c32f77a80_0 .net "in_a", 0 0, L_0x5c7c33140c90;  alias, 1 drivers
v0x5c7c32f77b70_0 .net "in_b", 0 0, L_0x5c7c33140c90;  alias, 1 drivers
v0x5c7c32f77c60_0 .net "out", 0 0, L_0x5c7c33140d40;  alias, 1 drivers
S_0x5c7c32f78300 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f76c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f79330_0 .net "in_a", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
v0x5c7c32f793d0_0 .net "in_b", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
v0x5c7c32f79490_0 .net "out", 0 0, L_0x5c7c33141060;  alias, 1 drivers
v0x5c7c32f795b0_0 .net "temp_out", 0 0, L_0x5c7c33140fb0;  1 drivers
S_0x5c7c32f784e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f78300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140fb0 .functor NAND 1, L_0x5c7c33140be0, L_0x5c7c33140be0, C4<1>, C4<1>;
v0x5c7c32f78750_0 .net "in_a", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
v0x5c7c32f78810_0 .net "in_b", 0 0, L_0x5c7c33140be0;  alias, 1 drivers
v0x5c7c32f78960_0 .net "out", 0 0, L_0x5c7c33140fb0;  alias, 1 drivers
S_0x5c7c32f78a60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f78300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f79180_0 .net "in_a", 0 0, L_0x5c7c33140fb0;  alias, 1 drivers
v0x5c7c32f79220_0 .net "out", 0 0, L_0x5c7c33141060;  alias, 1 drivers
S_0x5c7c32f78c30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f78a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141060 .functor NAND 1, L_0x5c7c33140fb0, L_0x5c7c33140fb0, C4<1>, C4<1>;
v0x5c7c32f78ea0_0 .net "in_a", 0 0, L_0x5c7c33140fb0;  alias, 1 drivers
v0x5c7c32f78f90_0 .net "in_b", 0 0, L_0x5c7c33140fb0;  alias, 1 drivers
v0x5c7c32f79080_0 .net "out", 0 0, L_0x5c7c33141060;  alias, 1 drivers
S_0x5c7c32f79720 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f76c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f7a760_0 .net "in_a", 0 0, L_0x5c7c33140df0;  alias, 1 drivers
v0x5c7c32f7a830_0 .net "in_b", 0 0, L_0x5c7c33141110;  alias, 1 drivers
v0x5c7c32f7a900_0 .net "out", 0 0, L_0x5c7c33141380;  alias, 1 drivers
v0x5c7c32f7aa20_0 .net "temp_out", 0 0, L_0x5c7c331412d0;  1 drivers
S_0x5c7c32f79900 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f79720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331412d0 .functor NAND 1, L_0x5c7c33140df0, L_0x5c7c33141110, C4<1>, C4<1>;
v0x5c7c32f79b50_0 .net "in_a", 0 0, L_0x5c7c33140df0;  alias, 1 drivers
v0x5c7c32f79c30_0 .net "in_b", 0 0, L_0x5c7c33141110;  alias, 1 drivers
v0x5c7c32f79cf0_0 .net "out", 0 0, L_0x5c7c331412d0;  alias, 1 drivers
S_0x5c7c32f79e40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f79720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f7a5b0_0 .net "in_a", 0 0, L_0x5c7c331412d0;  alias, 1 drivers
v0x5c7c32f7a650_0 .net "out", 0 0, L_0x5c7c33141380;  alias, 1 drivers
S_0x5c7c32f7a060 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f79e40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141380 .functor NAND 1, L_0x5c7c331412d0, L_0x5c7c331412d0, C4<1>, C4<1>;
v0x5c7c32f7a2d0_0 .net "in_a", 0 0, L_0x5c7c331412d0;  alias, 1 drivers
v0x5c7c32f7a3c0_0 .net "in_b", 0 0, L_0x5c7c331412d0;  alias, 1 drivers
v0x5c7c32f7a4b0_0 .net "out", 0 0, L_0x5c7c33141380;  alias, 1 drivers
S_0x5c7c32f7ab70 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f76c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f7b2a0_0 .net "in_a", 0 0, L_0x5c7c33140d40;  alias, 1 drivers
v0x5c7c32f7b340_0 .net "out", 0 0, L_0x5c7c33140df0;  alias, 1 drivers
S_0x5c7c32f7ad40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f7ab70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33140df0 .functor NAND 1, L_0x5c7c33140d40, L_0x5c7c33140d40, C4<1>, C4<1>;
v0x5c7c32f7afb0_0 .net "in_a", 0 0, L_0x5c7c33140d40;  alias, 1 drivers
v0x5c7c32f7b070_0 .net "in_b", 0 0, L_0x5c7c33140d40;  alias, 1 drivers
v0x5c7c32f7b1c0_0 .net "out", 0 0, L_0x5c7c33140df0;  alias, 1 drivers
S_0x5c7c32f7b440 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f76c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f7bc10_0 .net "in_a", 0 0, L_0x5c7c33141060;  alias, 1 drivers
v0x5c7c32f7bcb0_0 .net "out", 0 0, L_0x5c7c33141110;  alias, 1 drivers
S_0x5c7c32f7b6b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f7b440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141110 .functor NAND 1, L_0x5c7c33141060, L_0x5c7c33141060, C4<1>, C4<1>;
v0x5c7c32f7b920_0 .net "in_a", 0 0, L_0x5c7c33141060;  alias, 1 drivers
v0x5c7c32f7b9e0_0 .net "in_b", 0 0, L_0x5c7c33141060;  alias, 1 drivers
v0x5c7c32f7bb30_0 .net "out", 0 0, L_0x5c7c33141110;  alias, 1 drivers
S_0x5c7c32f7bdb0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f76c20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f7c550_0 .net "in_a", 0 0, L_0x5c7c33141380;  alias, 1 drivers
v0x5c7c32f7c5f0_0 .net "out", 0 0, L_0x5c7c33141430;  alias, 1 drivers
S_0x5c7c32f7bfd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f7bdb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141430 .functor NAND 1, L_0x5c7c33141380, L_0x5c7c33141380, C4<1>, C4<1>;
v0x5c7c32f7c240_0 .net "in_a", 0 0, L_0x5c7c33141380;  alias, 1 drivers
v0x5c7c32f7c300_0 .net "in_b", 0 0, L_0x5c7c33141380;  alias, 1 drivers
v0x5c7c32f7c450_0 .net "out", 0 0, L_0x5c7c33141430;  alias, 1 drivers
S_0x5c7c32f7d590 .scope module, "mux_gate4" "Mux" 15 11, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f87100_0 .net "in_a", 0 0, L_0x5c7c33142400;  1 drivers
v0x5c7c32f871a0_0 .net "in_b", 0 0, L_0x5c7c331424a0;  1 drivers
v0x5c7c32f872b0_0 .net "out", 0 0, L_0x5c7c33142240;  1 drivers
v0x5c7c32f87350_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f873f0_0 .net "sel_out", 0 0, L_0x5c7c33141730;  1 drivers
v0x5c7c32f87570_0 .net "temp_a_out", 0 0, L_0x5c7c33141890;  1 drivers
v0x5c7c32f87720_0 .net "temp_b_out", 0 0, L_0x5c7c331419f0;  1 drivers
S_0x5c7c32f7d790 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f7d590;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f7e7f0_0 .net "in_a", 0 0, L_0x5c7c33142400;  alias, 1 drivers
v0x5c7c32f7e8c0_0 .net "in_b", 0 0, L_0x5c7c33141730;  alias, 1 drivers
v0x5c7c32f7e990_0 .net "out", 0 0, L_0x5c7c33141890;  alias, 1 drivers
v0x5c7c32f7eab0_0 .net "temp_out", 0 0, L_0x5c7c331417e0;  1 drivers
S_0x5c7c32f7da00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f7d790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331417e0 .functor NAND 1, L_0x5c7c33142400, L_0x5c7c33141730, C4<1>, C4<1>;
v0x5c7c32f7dc70_0 .net "in_a", 0 0, L_0x5c7c33142400;  alias, 1 drivers
v0x5c7c32f7dd50_0 .net "in_b", 0 0, L_0x5c7c33141730;  alias, 1 drivers
v0x5c7c32f7de10_0 .net "out", 0 0, L_0x5c7c331417e0;  alias, 1 drivers
S_0x5c7c32f7df30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f7d790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f7e670_0 .net "in_a", 0 0, L_0x5c7c331417e0;  alias, 1 drivers
v0x5c7c32f7e710_0 .net "out", 0 0, L_0x5c7c33141890;  alias, 1 drivers
S_0x5c7c32f7e150 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f7df30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141890 .functor NAND 1, L_0x5c7c331417e0, L_0x5c7c331417e0, C4<1>, C4<1>;
v0x5c7c32f7e3c0_0 .net "in_a", 0 0, L_0x5c7c331417e0;  alias, 1 drivers
v0x5c7c32f7e480_0 .net "in_b", 0 0, L_0x5c7c331417e0;  alias, 1 drivers
v0x5c7c32f7e570_0 .net "out", 0 0, L_0x5c7c33141890;  alias, 1 drivers
S_0x5c7c32f7eb70 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f7d590;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f7fb80_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f7fc20_0 .net "in_b", 0 0, L_0x5c7c331424a0;  alias, 1 drivers
v0x5c7c32f7fd10_0 .net "out", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
v0x5c7c32f7fe30_0 .net "temp_out", 0 0, L_0x5c7c33141940;  1 drivers
S_0x5c7c32f7ed50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f7eb70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141940 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c331424a0, C4<1>, C4<1>;
v0x5c7c32f7efc0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f7f080_0 .net "in_b", 0 0, L_0x5c7c331424a0;  alias, 1 drivers
v0x5c7c32f7f140_0 .net "out", 0 0, L_0x5c7c33141940;  alias, 1 drivers
S_0x5c7c32f7f260 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f7eb70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f7f9d0_0 .net "in_a", 0 0, L_0x5c7c33141940;  alias, 1 drivers
v0x5c7c32f7fa70_0 .net "out", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
S_0x5c7c32f7f480 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f7f260;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331419f0 .functor NAND 1, L_0x5c7c33141940, L_0x5c7c33141940, C4<1>, C4<1>;
v0x5c7c32f7f6f0_0 .net "in_a", 0 0, L_0x5c7c33141940;  alias, 1 drivers
v0x5c7c32f7f7e0_0 .net "in_b", 0 0, L_0x5c7c33141940;  alias, 1 drivers
v0x5c7c32f7f8d0_0 .net "out", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
S_0x5c7c32f7fef0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f7d590;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f805f0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f80ea0_0 .net "out", 0 0, L_0x5c7c33141730;  alias, 1 drivers
S_0x5c7c32f800c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f7fef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141730 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f80310_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f803d0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f80490_0 .net "out", 0 0, L_0x5c7c33141730;  alias, 1 drivers
S_0x5c7c32f80fa0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f7d590;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f86a50_0 .net "branch1_out", 0 0, L_0x5c7c33141c00;  1 drivers
v0x5c7c32f86b80_0 .net "branch2_out", 0 0, L_0x5c7c33141f20;  1 drivers
v0x5c7c32f86cd0_0 .net "in_a", 0 0, L_0x5c7c33141890;  alias, 1 drivers
v0x5c7c32f86da0_0 .net "in_b", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
v0x5c7c32f86e40_0 .net "out", 0 0, L_0x5c7c33142240;  alias, 1 drivers
v0x5c7c32f86ee0_0 .net "temp1_out", 0 0, L_0x5c7c33141b50;  1 drivers
v0x5c7c32f86f80_0 .net "temp2_out", 0 0, L_0x5c7c33141e70;  1 drivers
v0x5c7c32f87020_0 .net "temp3_out", 0 0, L_0x5c7c33142190;  1 drivers
S_0x5c7c32f811d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f80fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f82290_0 .net "in_a", 0 0, L_0x5c7c33141890;  alias, 1 drivers
v0x5c7c32f82330_0 .net "in_b", 0 0, L_0x5c7c33141890;  alias, 1 drivers
v0x5c7c32f823f0_0 .net "out", 0 0, L_0x5c7c33141b50;  alias, 1 drivers
v0x5c7c32f82510_0 .net "temp_out", 0 0, L_0x5c7c33141aa0;  1 drivers
S_0x5c7c32f81440 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f811d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141aa0 .functor NAND 1, L_0x5c7c33141890, L_0x5c7c33141890, C4<1>, C4<1>;
v0x5c7c32f816b0_0 .net "in_a", 0 0, L_0x5c7c33141890;  alias, 1 drivers
v0x5c7c32f81770_0 .net "in_b", 0 0, L_0x5c7c33141890;  alias, 1 drivers
v0x5c7c32f818c0_0 .net "out", 0 0, L_0x5c7c33141aa0;  alias, 1 drivers
S_0x5c7c32f819c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f811d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f820e0_0 .net "in_a", 0 0, L_0x5c7c33141aa0;  alias, 1 drivers
v0x5c7c32f82180_0 .net "out", 0 0, L_0x5c7c33141b50;  alias, 1 drivers
S_0x5c7c32f81b90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f819c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141b50 .functor NAND 1, L_0x5c7c33141aa0, L_0x5c7c33141aa0, C4<1>, C4<1>;
v0x5c7c32f81e00_0 .net "in_a", 0 0, L_0x5c7c33141aa0;  alias, 1 drivers
v0x5c7c32f81ef0_0 .net "in_b", 0 0, L_0x5c7c33141aa0;  alias, 1 drivers
v0x5c7c32f81fe0_0 .net "out", 0 0, L_0x5c7c33141b50;  alias, 1 drivers
S_0x5c7c32f82680 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f80fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f836b0_0 .net "in_a", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
v0x5c7c32f83750_0 .net "in_b", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
v0x5c7c32f83810_0 .net "out", 0 0, L_0x5c7c33141e70;  alias, 1 drivers
v0x5c7c32f83930_0 .net "temp_out", 0 0, L_0x5c7c33141dc0;  1 drivers
S_0x5c7c32f82860 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f82680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141dc0 .functor NAND 1, L_0x5c7c331419f0, L_0x5c7c331419f0, C4<1>, C4<1>;
v0x5c7c32f82ad0_0 .net "in_a", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
v0x5c7c32f82b90_0 .net "in_b", 0 0, L_0x5c7c331419f0;  alias, 1 drivers
v0x5c7c32f82ce0_0 .net "out", 0 0, L_0x5c7c33141dc0;  alias, 1 drivers
S_0x5c7c32f82de0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f82680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f83500_0 .net "in_a", 0 0, L_0x5c7c33141dc0;  alias, 1 drivers
v0x5c7c32f835a0_0 .net "out", 0 0, L_0x5c7c33141e70;  alias, 1 drivers
S_0x5c7c32f82fb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f82de0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141e70 .functor NAND 1, L_0x5c7c33141dc0, L_0x5c7c33141dc0, C4<1>, C4<1>;
v0x5c7c32f83220_0 .net "in_a", 0 0, L_0x5c7c33141dc0;  alias, 1 drivers
v0x5c7c32f83310_0 .net "in_b", 0 0, L_0x5c7c33141dc0;  alias, 1 drivers
v0x5c7c32f83400_0 .net "out", 0 0, L_0x5c7c33141e70;  alias, 1 drivers
S_0x5c7c32f83aa0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f80fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f84ae0_0 .net "in_a", 0 0, L_0x5c7c33141c00;  alias, 1 drivers
v0x5c7c32f84bb0_0 .net "in_b", 0 0, L_0x5c7c33141f20;  alias, 1 drivers
v0x5c7c32f84c80_0 .net "out", 0 0, L_0x5c7c33142190;  alias, 1 drivers
v0x5c7c32f84da0_0 .net "temp_out", 0 0, L_0x5c7c331420e0;  1 drivers
S_0x5c7c32f83c80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f83aa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331420e0 .functor NAND 1, L_0x5c7c33141c00, L_0x5c7c33141f20, C4<1>, C4<1>;
v0x5c7c32f83ed0_0 .net "in_a", 0 0, L_0x5c7c33141c00;  alias, 1 drivers
v0x5c7c32f83fb0_0 .net "in_b", 0 0, L_0x5c7c33141f20;  alias, 1 drivers
v0x5c7c32f84070_0 .net "out", 0 0, L_0x5c7c331420e0;  alias, 1 drivers
S_0x5c7c32f841c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f83aa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f84930_0 .net "in_a", 0 0, L_0x5c7c331420e0;  alias, 1 drivers
v0x5c7c32f849d0_0 .net "out", 0 0, L_0x5c7c33142190;  alias, 1 drivers
S_0x5c7c32f843e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f841c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142190 .functor NAND 1, L_0x5c7c331420e0, L_0x5c7c331420e0, C4<1>, C4<1>;
v0x5c7c32f84650_0 .net "in_a", 0 0, L_0x5c7c331420e0;  alias, 1 drivers
v0x5c7c32f84740_0 .net "in_b", 0 0, L_0x5c7c331420e0;  alias, 1 drivers
v0x5c7c32f84830_0 .net "out", 0 0, L_0x5c7c33142190;  alias, 1 drivers
S_0x5c7c32f84ef0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f80fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f85620_0 .net "in_a", 0 0, L_0x5c7c33141b50;  alias, 1 drivers
v0x5c7c32f856c0_0 .net "out", 0 0, L_0x5c7c33141c00;  alias, 1 drivers
S_0x5c7c32f850c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f84ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141c00 .functor NAND 1, L_0x5c7c33141b50, L_0x5c7c33141b50, C4<1>, C4<1>;
v0x5c7c32f85330_0 .net "in_a", 0 0, L_0x5c7c33141b50;  alias, 1 drivers
v0x5c7c32f853f0_0 .net "in_b", 0 0, L_0x5c7c33141b50;  alias, 1 drivers
v0x5c7c32f85540_0 .net "out", 0 0, L_0x5c7c33141c00;  alias, 1 drivers
S_0x5c7c32f857c0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f80fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f85f90_0 .net "in_a", 0 0, L_0x5c7c33141e70;  alias, 1 drivers
v0x5c7c32f86030_0 .net "out", 0 0, L_0x5c7c33141f20;  alias, 1 drivers
S_0x5c7c32f85a30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f857c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33141f20 .functor NAND 1, L_0x5c7c33141e70, L_0x5c7c33141e70, C4<1>, C4<1>;
v0x5c7c32f85ca0_0 .net "in_a", 0 0, L_0x5c7c33141e70;  alias, 1 drivers
v0x5c7c32f85d60_0 .net "in_b", 0 0, L_0x5c7c33141e70;  alias, 1 drivers
v0x5c7c32f85eb0_0 .net "out", 0 0, L_0x5c7c33141f20;  alias, 1 drivers
S_0x5c7c32f86130 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f80fa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f868d0_0 .net "in_a", 0 0, L_0x5c7c33142190;  alias, 1 drivers
v0x5c7c32f86970_0 .net "out", 0 0, L_0x5c7c33142240;  alias, 1 drivers
S_0x5c7c32f86350 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f86130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142240 .functor NAND 1, L_0x5c7c33142190, L_0x5c7c33142190, C4<1>, C4<1>;
v0x5c7c32f865c0_0 .net "in_a", 0 0, L_0x5c7c33142190;  alias, 1 drivers
v0x5c7c32f86680_0 .net "in_b", 0 0, L_0x5c7c33142190;  alias, 1 drivers
v0x5c7c32f867d0_0 .net "out", 0 0, L_0x5c7c33142240;  alias, 1 drivers
S_0x5c7c32f87910 .scope module, "mux_gate5" "Mux" 15 12, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f90c70_0 .net "in_a", 0 0, L_0x5c7c33143270;  1 drivers
v0x5c7c32f90d10_0 .net "in_b", 0 0, L_0x5c7c33143310;  1 drivers
v0x5c7c32f90e20_0 .net "out", 0 0, L_0x5c7c331430b0;  1 drivers
v0x5c7c32f90ec0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f90f60_0 .net "sel_out", 0 0, L_0x5c7c331425a0;  1 drivers
v0x5c7c32f910e0_0 .net "temp_a_out", 0 0, L_0x5c7c33142700;  1 drivers
v0x5c7c32f91290_0 .net "temp_b_out", 0 0, L_0x5c7c33142860;  1 drivers
S_0x5c7c32f87b10 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f87910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f88b70_0 .net "in_a", 0 0, L_0x5c7c33143270;  alias, 1 drivers
v0x5c7c32f88c40_0 .net "in_b", 0 0, L_0x5c7c331425a0;  alias, 1 drivers
v0x5c7c32f88d10_0 .net "out", 0 0, L_0x5c7c33142700;  alias, 1 drivers
v0x5c7c32f88e30_0 .net "temp_out", 0 0, L_0x5c7c33142650;  1 drivers
S_0x5c7c32f87d80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f87b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142650 .functor NAND 1, L_0x5c7c33143270, L_0x5c7c331425a0, C4<1>, C4<1>;
v0x5c7c32f87ff0_0 .net "in_a", 0 0, L_0x5c7c33143270;  alias, 1 drivers
v0x5c7c32f880d0_0 .net "in_b", 0 0, L_0x5c7c331425a0;  alias, 1 drivers
v0x5c7c32f88190_0 .net "out", 0 0, L_0x5c7c33142650;  alias, 1 drivers
S_0x5c7c32f882b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f87b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f889f0_0 .net "in_a", 0 0, L_0x5c7c33142650;  alias, 1 drivers
v0x5c7c32f88a90_0 .net "out", 0 0, L_0x5c7c33142700;  alias, 1 drivers
S_0x5c7c32f884d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f882b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142700 .functor NAND 1, L_0x5c7c33142650, L_0x5c7c33142650, C4<1>, C4<1>;
v0x5c7c32f88740_0 .net "in_a", 0 0, L_0x5c7c33142650;  alias, 1 drivers
v0x5c7c32f88800_0 .net "in_b", 0 0, L_0x5c7c33142650;  alias, 1 drivers
v0x5c7c32f888f0_0 .net "out", 0 0, L_0x5c7c33142700;  alias, 1 drivers
S_0x5c7c32f88ef0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f87910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f89f00_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f89fa0_0 .net "in_b", 0 0, L_0x5c7c33143310;  alias, 1 drivers
v0x5c7c32f8a090_0 .net "out", 0 0, L_0x5c7c33142860;  alias, 1 drivers
v0x5c7c32f8a1b0_0 .net "temp_out", 0 0, L_0x5c7c331427b0;  1 drivers
S_0x5c7c32f890d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f88ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331427b0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33143310, C4<1>, C4<1>;
v0x5c7c32f89340_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f89400_0 .net "in_b", 0 0, L_0x5c7c33143310;  alias, 1 drivers
v0x5c7c32f894c0_0 .net "out", 0 0, L_0x5c7c331427b0;  alias, 1 drivers
S_0x5c7c32f895e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f88ef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f89d50_0 .net "in_a", 0 0, L_0x5c7c331427b0;  alias, 1 drivers
v0x5c7c32f89df0_0 .net "out", 0 0, L_0x5c7c33142860;  alias, 1 drivers
S_0x5c7c32f89800 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f895e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142860 .functor NAND 1, L_0x5c7c331427b0, L_0x5c7c331427b0, C4<1>, C4<1>;
v0x5c7c32f89a70_0 .net "in_a", 0 0, L_0x5c7c331427b0;  alias, 1 drivers
v0x5c7c32f89b60_0 .net "in_b", 0 0, L_0x5c7c331427b0;  alias, 1 drivers
v0x5c7c32f89c50_0 .net "out", 0 0, L_0x5c7c33142860;  alias, 1 drivers
S_0x5c7c32f8a270 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f87910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f8a970_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f8aa10_0 .net "out", 0 0, L_0x5c7c331425a0;  alias, 1 drivers
S_0x5c7c32f8a440 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8a270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331425a0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f8a690_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f8a750_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f8a810_0 .net "out", 0 0, L_0x5c7c331425a0;  alias, 1 drivers
S_0x5c7c32f8ab10 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f87910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f905c0_0 .net "branch1_out", 0 0, L_0x5c7c33142a70;  1 drivers
v0x5c7c32f906f0_0 .net "branch2_out", 0 0, L_0x5c7c33142d90;  1 drivers
v0x5c7c32f90840_0 .net "in_a", 0 0, L_0x5c7c33142700;  alias, 1 drivers
v0x5c7c32f90910_0 .net "in_b", 0 0, L_0x5c7c33142860;  alias, 1 drivers
v0x5c7c32f909b0_0 .net "out", 0 0, L_0x5c7c331430b0;  alias, 1 drivers
v0x5c7c32f90a50_0 .net "temp1_out", 0 0, L_0x5c7c331429c0;  1 drivers
v0x5c7c32f90af0_0 .net "temp2_out", 0 0, L_0x5c7c33142ce0;  1 drivers
v0x5c7c32f90b90_0 .net "temp3_out", 0 0, L_0x5c7c33143000;  1 drivers
S_0x5c7c32f8ad40 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f8ab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f8be00_0 .net "in_a", 0 0, L_0x5c7c33142700;  alias, 1 drivers
v0x5c7c32f8bea0_0 .net "in_b", 0 0, L_0x5c7c33142700;  alias, 1 drivers
v0x5c7c32f8bf60_0 .net "out", 0 0, L_0x5c7c331429c0;  alias, 1 drivers
v0x5c7c32f8c080_0 .net "temp_out", 0 0, L_0x5c7c33142910;  1 drivers
S_0x5c7c32f8afb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f8ad40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142910 .functor NAND 1, L_0x5c7c33142700, L_0x5c7c33142700, C4<1>, C4<1>;
v0x5c7c32f8b220_0 .net "in_a", 0 0, L_0x5c7c33142700;  alias, 1 drivers
v0x5c7c32f8b2e0_0 .net "in_b", 0 0, L_0x5c7c33142700;  alias, 1 drivers
v0x5c7c32f8b430_0 .net "out", 0 0, L_0x5c7c33142910;  alias, 1 drivers
S_0x5c7c32f8b530 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f8ad40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f8bc50_0 .net "in_a", 0 0, L_0x5c7c33142910;  alias, 1 drivers
v0x5c7c32f8bcf0_0 .net "out", 0 0, L_0x5c7c331429c0;  alias, 1 drivers
S_0x5c7c32f8b700 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8b530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331429c0 .functor NAND 1, L_0x5c7c33142910, L_0x5c7c33142910, C4<1>, C4<1>;
v0x5c7c32f8b970_0 .net "in_a", 0 0, L_0x5c7c33142910;  alias, 1 drivers
v0x5c7c32f8ba60_0 .net "in_b", 0 0, L_0x5c7c33142910;  alias, 1 drivers
v0x5c7c32f8bb50_0 .net "out", 0 0, L_0x5c7c331429c0;  alias, 1 drivers
S_0x5c7c32f8c1f0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f8ab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f8d220_0 .net "in_a", 0 0, L_0x5c7c33142860;  alias, 1 drivers
v0x5c7c32f8d2c0_0 .net "in_b", 0 0, L_0x5c7c33142860;  alias, 1 drivers
v0x5c7c32f8d380_0 .net "out", 0 0, L_0x5c7c33142ce0;  alias, 1 drivers
v0x5c7c32f8d4a0_0 .net "temp_out", 0 0, L_0x5c7c33142c30;  1 drivers
S_0x5c7c32f8c3d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f8c1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142c30 .functor NAND 1, L_0x5c7c33142860, L_0x5c7c33142860, C4<1>, C4<1>;
v0x5c7c32f8c640_0 .net "in_a", 0 0, L_0x5c7c33142860;  alias, 1 drivers
v0x5c7c32f8c700_0 .net "in_b", 0 0, L_0x5c7c33142860;  alias, 1 drivers
v0x5c7c32f8c850_0 .net "out", 0 0, L_0x5c7c33142c30;  alias, 1 drivers
S_0x5c7c32f8c950 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f8c1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f8d070_0 .net "in_a", 0 0, L_0x5c7c33142c30;  alias, 1 drivers
v0x5c7c32f8d110_0 .net "out", 0 0, L_0x5c7c33142ce0;  alias, 1 drivers
S_0x5c7c32f8cb20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8c950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142ce0 .functor NAND 1, L_0x5c7c33142c30, L_0x5c7c33142c30, C4<1>, C4<1>;
v0x5c7c32f8cd90_0 .net "in_a", 0 0, L_0x5c7c33142c30;  alias, 1 drivers
v0x5c7c32f8ce80_0 .net "in_b", 0 0, L_0x5c7c33142c30;  alias, 1 drivers
v0x5c7c32f8cf70_0 .net "out", 0 0, L_0x5c7c33142ce0;  alias, 1 drivers
S_0x5c7c32f8d610 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f8ab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f8e650_0 .net "in_a", 0 0, L_0x5c7c33142a70;  alias, 1 drivers
v0x5c7c32f8e720_0 .net "in_b", 0 0, L_0x5c7c33142d90;  alias, 1 drivers
v0x5c7c32f8e7f0_0 .net "out", 0 0, L_0x5c7c33143000;  alias, 1 drivers
v0x5c7c32f8e910_0 .net "temp_out", 0 0, L_0x5c7c33142f50;  1 drivers
S_0x5c7c32f8d7f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f8d610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142f50 .functor NAND 1, L_0x5c7c33142a70, L_0x5c7c33142d90, C4<1>, C4<1>;
v0x5c7c32f8da40_0 .net "in_a", 0 0, L_0x5c7c33142a70;  alias, 1 drivers
v0x5c7c32f8db20_0 .net "in_b", 0 0, L_0x5c7c33142d90;  alias, 1 drivers
v0x5c7c32f8dbe0_0 .net "out", 0 0, L_0x5c7c33142f50;  alias, 1 drivers
S_0x5c7c32f8dd30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f8d610;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f8e4a0_0 .net "in_a", 0 0, L_0x5c7c33142f50;  alias, 1 drivers
v0x5c7c32f8e540_0 .net "out", 0 0, L_0x5c7c33143000;  alias, 1 drivers
S_0x5c7c32f8df50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8dd30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143000 .functor NAND 1, L_0x5c7c33142f50, L_0x5c7c33142f50, C4<1>, C4<1>;
v0x5c7c32f8e1c0_0 .net "in_a", 0 0, L_0x5c7c33142f50;  alias, 1 drivers
v0x5c7c32f8e2b0_0 .net "in_b", 0 0, L_0x5c7c33142f50;  alias, 1 drivers
v0x5c7c32f8e3a0_0 .net "out", 0 0, L_0x5c7c33143000;  alias, 1 drivers
S_0x5c7c32f8ea60 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f8ab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f8f190_0 .net "in_a", 0 0, L_0x5c7c331429c0;  alias, 1 drivers
v0x5c7c32f8f230_0 .net "out", 0 0, L_0x5c7c33142a70;  alias, 1 drivers
S_0x5c7c32f8ec30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8ea60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142a70 .functor NAND 1, L_0x5c7c331429c0, L_0x5c7c331429c0, C4<1>, C4<1>;
v0x5c7c32f8eea0_0 .net "in_a", 0 0, L_0x5c7c331429c0;  alias, 1 drivers
v0x5c7c32f8ef60_0 .net "in_b", 0 0, L_0x5c7c331429c0;  alias, 1 drivers
v0x5c7c32f8f0b0_0 .net "out", 0 0, L_0x5c7c33142a70;  alias, 1 drivers
S_0x5c7c32f8f330 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f8ab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f8fb00_0 .net "in_a", 0 0, L_0x5c7c33142ce0;  alias, 1 drivers
v0x5c7c32f8fba0_0 .net "out", 0 0, L_0x5c7c33142d90;  alias, 1 drivers
S_0x5c7c32f8f5a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8f330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33142d90 .functor NAND 1, L_0x5c7c33142ce0, L_0x5c7c33142ce0, C4<1>, C4<1>;
v0x5c7c32f8f810_0 .net "in_a", 0 0, L_0x5c7c33142ce0;  alias, 1 drivers
v0x5c7c32f8f8d0_0 .net "in_b", 0 0, L_0x5c7c33142ce0;  alias, 1 drivers
v0x5c7c32f8fa20_0 .net "out", 0 0, L_0x5c7c33142d90;  alias, 1 drivers
S_0x5c7c32f8fca0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f8ab10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f90440_0 .net "in_a", 0 0, L_0x5c7c33143000;  alias, 1 drivers
v0x5c7c32f904e0_0 .net "out", 0 0, L_0x5c7c331430b0;  alias, 1 drivers
S_0x5c7c32f8fec0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f8fca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331430b0 .functor NAND 1, L_0x5c7c33143000, L_0x5c7c33143000, C4<1>, C4<1>;
v0x5c7c32f90130_0 .net "in_a", 0 0, L_0x5c7c33143000;  alias, 1 drivers
v0x5c7c32f901f0_0 .net "in_b", 0 0, L_0x5c7c33143000;  alias, 1 drivers
v0x5c7c32f90340_0 .net "out", 0 0, L_0x5c7c331430b0;  alias, 1 drivers
S_0x5c7c32f91480 .scope module, "mux_gate6" "Mux" 15 13, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32f9a7e0_0 .net "in_a", 0 0, L_0x5c7c331440f0;  1 drivers
v0x5c7c32f9a880_0 .net "in_b", 0 0, L_0x5c7c331442a0;  1 drivers
v0x5c7c32f9a990_0 .net "out", 0 0, L_0x5c7c33143f30;  1 drivers
v0x5c7c32f9aa30_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f9aad0_0 .net "sel_out", 0 0, L_0x5c7c33143420;  1 drivers
v0x5c7c32f9ac50_0 .net "temp_a_out", 0 0, L_0x5c7c33143580;  1 drivers
v0x5c7c32f9ae00_0 .net "temp_b_out", 0 0, L_0x5c7c331436e0;  1 drivers
S_0x5c7c32f91680 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f91480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f926e0_0 .net "in_a", 0 0, L_0x5c7c331440f0;  alias, 1 drivers
v0x5c7c32f927b0_0 .net "in_b", 0 0, L_0x5c7c33143420;  alias, 1 drivers
v0x5c7c32f92880_0 .net "out", 0 0, L_0x5c7c33143580;  alias, 1 drivers
v0x5c7c32f929a0_0 .net "temp_out", 0 0, L_0x5c7c331434d0;  1 drivers
S_0x5c7c32f918f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f91680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331434d0 .functor NAND 1, L_0x5c7c331440f0, L_0x5c7c33143420, C4<1>, C4<1>;
v0x5c7c32f91b60_0 .net "in_a", 0 0, L_0x5c7c331440f0;  alias, 1 drivers
v0x5c7c32f91c40_0 .net "in_b", 0 0, L_0x5c7c33143420;  alias, 1 drivers
v0x5c7c32f91d00_0 .net "out", 0 0, L_0x5c7c331434d0;  alias, 1 drivers
S_0x5c7c32f91e20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f91680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f92560_0 .net "in_a", 0 0, L_0x5c7c331434d0;  alias, 1 drivers
v0x5c7c32f92600_0 .net "out", 0 0, L_0x5c7c33143580;  alias, 1 drivers
S_0x5c7c32f92040 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f91e20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143580 .functor NAND 1, L_0x5c7c331434d0, L_0x5c7c331434d0, C4<1>, C4<1>;
v0x5c7c32f922b0_0 .net "in_a", 0 0, L_0x5c7c331434d0;  alias, 1 drivers
v0x5c7c32f92370_0 .net "in_b", 0 0, L_0x5c7c331434d0;  alias, 1 drivers
v0x5c7c32f92460_0 .net "out", 0 0, L_0x5c7c33143580;  alias, 1 drivers
S_0x5c7c32f92a60 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f91480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f93a70_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f93b10_0 .net "in_b", 0 0, L_0x5c7c331442a0;  alias, 1 drivers
v0x5c7c32f93c00_0 .net "out", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
v0x5c7c32f93d20_0 .net "temp_out", 0 0, L_0x5c7c33143630;  1 drivers
S_0x5c7c32f92c40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f92a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143630 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c331442a0, C4<1>, C4<1>;
v0x5c7c32f92eb0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f92f70_0 .net "in_b", 0 0, L_0x5c7c331442a0;  alias, 1 drivers
v0x5c7c32f93030_0 .net "out", 0 0, L_0x5c7c33143630;  alias, 1 drivers
S_0x5c7c32f93150 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f92a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f938c0_0 .net "in_a", 0 0, L_0x5c7c33143630;  alias, 1 drivers
v0x5c7c32f93960_0 .net "out", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
S_0x5c7c32f93370 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f93150;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331436e0 .functor NAND 1, L_0x5c7c33143630, L_0x5c7c33143630, C4<1>, C4<1>;
v0x5c7c32f935e0_0 .net "in_a", 0 0, L_0x5c7c33143630;  alias, 1 drivers
v0x5c7c32f936d0_0 .net "in_b", 0 0, L_0x5c7c33143630;  alias, 1 drivers
v0x5c7c32f937c0_0 .net "out", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
S_0x5c7c32f93de0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f91480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f944e0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f94580_0 .net "out", 0 0, L_0x5c7c33143420;  alias, 1 drivers
S_0x5c7c32f93fb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f93de0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143420 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f94200_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f942c0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f94380_0 .net "out", 0 0, L_0x5c7c33143420;  alias, 1 drivers
S_0x5c7c32f94680 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f91480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f9a130_0 .net "branch1_out", 0 0, L_0x5c7c331438f0;  1 drivers
v0x5c7c32f9a260_0 .net "branch2_out", 0 0, L_0x5c7c33143c10;  1 drivers
v0x5c7c32f9a3b0_0 .net "in_a", 0 0, L_0x5c7c33143580;  alias, 1 drivers
v0x5c7c32f9a480_0 .net "in_b", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
v0x5c7c32f9a520_0 .net "out", 0 0, L_0x5c7c33143f30;  alias, 1 drivers
v0x5c7c32f9a5c0_0 .net "temp1_out", 0 0, L_0x5c7c33143840;  1 drivers
v0x5c7c32f9a660_0 .net "temp2_out", 0 0, L_0x5c7c33143b60;  1 drivers
v0x5c7c32f9a700_0 .net "temp3_out", 0 0, L_0x5c7c33143e80;  1 drivers
S_0x5c7c32f948b0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f94680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f95970_0 .net "in_a", 0 0, L_0x5c7c33143580;  alias, 1 drivers
v0x5c7c32f95a10_0 .net "in_b", 0 0, L_0x5c7c33143580;  alias, 1 drivers
v0x5c7c32f95ad0_0 .net "out", 0 0, L_0x5c7c33143840;  alias, 1 drivers
v0x5c7c32f95bf0_0 .net "temp_out", 0 0, L_0x5c7c33143790;  1 drivers
S_0x5c7c32f94b20 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f948b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143790 .functor NAND 1, L_0x5c7c33143580, L_0x5c7c33143580, C4<1>, C4<1>;
v0x5c7c32f94d90_0 .net "in_a", 0 0, L_0x5c7c33143580;  alias, 1 drivers
v0x5c7c32f94e50_0 .net "in_b", 0 0, L_0x5c7c33143580;  alias, 1 drivers
v0x5c7c32f94fa0_0 .net "out", 0 0, L_0x5c7c33143790;  alias, 1 drivers
S_0x5c7c32f950a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f948b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f957c0_0 .net "in_a", 0 0, L_0x5c7c33143790;  alias, 1 drivers
v0x5c7c32f95860_0 .net "out", 0 0, L_0x5c7c33143840;  alias, 1 drivers
S_0x5c7c32f95270 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f950a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143840 .functor NAND 1, L_0x5c7c33143790, L_0x5c7c33143790, C4<1>, C4<1>;
v0x5c7c32f954e0_0 .net "in_a", 0 0, L_0x5c7c33143790;  alias, 1 drivers
v0x5c7c32f955d0_0 .net "in_b", 0 0, L_0x5c7c33143790;  alias, 1 drivers
v0x5c7c32f956c0_0 .net "out", 0 0, L_0x5c7c33143840;  alias, 1 drivers
S_0x5c7c32f95d60 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f94680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f96d90_0 .net "in_a", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
v0x5c7c32f96e30_0 .net "in_b", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
v0x5c7c32f96ef0_0 .net "out", 0 0, L_0x5c7c33143b60;  alias, 1 drivers
v0x5c7c32f97010_0 .net "temp_out", 0 0, L_0x5c7c33143ab0;  1 drivers
S_0x5c7c32f95f40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f95d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143ab0 .functor NAND 1, L_0x5c7c331436e0, L_0x5c7c331436e0, C4<1>, C4<1>;
v0x5c7c32f961b0_0 .net "in_a", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
v0x5c7c32f96270_0 .net "in_b", 0 0, L_0x5c7c331436e0;  alias, 1 drivers
v0x5c7c32f963c0_0 .net "out", 0 0, L_0x5c7c33143ab0;  alias, 1 drivers
S_0x5c7c32f964c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f95d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f96be0_0 .net "in_a", 0 0, L_0x5c7c33143ab0;  alias, 1 drivers
v0x5c7c32f96c80_0 .net "out", 0 0, L_0x5c7c33143b60;  alias, 1 drivers
S_0x5c7c32f96690 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f964c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143b60 .functor NAND 1, L_0x5c7c33143ab0, L_0x5c7c33143ab0, C4<1>, C4<1>;
v0x5c7c32f96900_0 .net "in_a", 0 0, L_0x5c7c33143ab0;  alias, 1 drivers
v0x5c7c32f969f0_0 .net "in_b", 0 0, L_0x5c7c33143ab0;  alias, 1 drivers
v0x5c7c32f96ae0_0 .net "out", 0 0, L_0x5c7c33143b60;  alias, 1 drivers
S_0x5c7c32f97180 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f94680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f981c0_0 .net "in_a", 0 0, L_0x5c7c331438f0;  alias, 1 drivers
v0x5c7c32f98290_0 .net "in_b", 0 0, L_0x5c7c33143c10;  alias, 1 drivers
v0x5c7c32f98360_0 .net "out", 0 0, L_0x5c7c33143e80;  alias, 1 drivers
v0x5c7c32f98480_0 .net "temp_out", 0 0, L_0x5c7c33143dd0;  1 drivers
S_0x5c7c32f97360 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f97180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143dd0 .functor NAND 1, L_0x5c7c331438f0, L_0x5c7c33143c10, C4<1>, C4<1>;
v0x5c7c32f975b0_0 .net "in_a", 0 0, L_0x5c7c331438f0;  alias, 1 drivers
v0x5c7c32f97690_0 .net "in_b", 0 0, L_0x5c7c33143c10;  alias, 1 drivers
v0x5c7c32f97750_0 .net "out", 0 0, L_0x5c7c33143dd0;  alias, 1 drivers
S_0x5c7c32f978a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f97180;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f98010_0 .net "in_a", 0 0, L_0x5c7c33143dd0;  alias, 1 drivers
v0x5c7c32f980b0_0 .net "out", 0 0, L_0x5c7c33143e80;  alias, 1 drivers
S_0x5c7c32f97ac0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f978a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143e80 .functor NAND 1, L_0x5c7c33143dd0, L_0x5c7c33143dd0, C4<1>, C4<1>;
v0x5c7c32f97d30_0 .net "in_a", 0 0, L_0x5c7c33143dd0;  alias, 1 drivers
v0x5c7c32f97e20_0 .net "in_b", 0 0, L_0x5c7c33143dd0;  alias, 1 drivers
v0x5c7c32f97f10_0 .net "out", 0 0, L_0x5c7c33143e80;  alias, 1 drivers
S_0x5c7c32f985d0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f94680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f98d00_0 .net "in_a", 0 0, L_0x5c7c33143840;  alias, 1 drivers
v0x5c7c32f98da0_0 .net "out", 0 0, L_0x5c7c331438f0;  alias, 1 drivers
S_0x5c7c32f987a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f985d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331438f0 .functor NAND 1, L_0x5c7c33143840, L_0x5c7c33143840, C4<1>, C4<1>;
v0x5c7c32f98a10_0 .net "in_a", 0 0, L_0x5c7c33143840;  alias, 1 drivers
v0x5c7c32f98ad0_0 .net "in_b", 0 0, L_0x5c7c33143840;  alias, 1 drivers
v0x5c7c32f98c20_0 .net "out", 0 0, L_0x5c7c331438f0;  alias, 1 drivers
S_0x5c7c32f98ea0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f94680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f99670_0 .net "in_a", 0 0, L_0x5c7c33143b60;  alias, 1 drivers
v0x5c7c32f99710_0 .net "out", 0 0, L_0x5c7c33143c10;  alias, 1 drivers
S_0x5c7c32f99110 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f98ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143c10 .functor NAND 1, L_0x5c7c33143b60, L_0x5c7c33143b60, C4<1>, C4<1>;
v0x5c7c32f99380_0 .net "in_a", 0 0, L_0x5c7c33143b60;  alias, 1 drivers
v0x5c7c32f99440_0 .net "in_b", 0 0, L_0x5c7c33143b60;  alias, 1 drivers
v0x5c7c32f99590_0 .net "out", 0 0, L_0x5c7c33143c10;  alias, 1 drivers
S_0x5c7c32f99810 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f94680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f99fb0_0 .net "in_a", 0 0, L_0x5c7c33143e80;  alias, 1 drivers
v0x5c7c32f9a050_0 .net "out", 0 0, L_0x5c7c33143f30;  alias, 1 drivers
S_0x5c7c32f99a30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f99810;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33143f30 .functor NAND 1, L_0x5c7c33143e80, L_0x5c7c33143e80, C4<1>, C4<1>;
v0x5c7c32f99ca0_0 .net "in_a", 0 0, L_0x5c7c33143e80;  alias, 1 drivers
v0x5c7c32f99d60_0 .net "in_b", 0 0, L_0x5c7c33143e80;  alias, 1 drivers
v0x5c7c32f99eb0_0 .net "out", 0 0, L_0x5c7c33143f30;  alias, 1 drivers
S_0x5c7c32f9aff0 .scope module, "mux_gate7" "Mux" 15 14, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fa4350_0 .net "in_a", 0 0, L_0x5c7c33145130;  1 drivers
v0x5c7c32fa43f0_0 .net "in_b", 0 0, L_0x5c7c331451d0;  1 drivers
v0x5c7c32fa4500_0 .net "out", 0 0, L_0x5c7c33144f70;  1 drivers
v0x5c7c32fa45a0_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fa4640_0 .net "sel_out", 0 0, L_0x5c7c331433b0;  1 drivers
v0x5c7c32fa47c0_0 .net "temp_a_out", 0 0, L_0x5c7c331445c0;  1 drivers
v0x5c7c32fa4970_0 .net "temp_b_out", 0 0, L_0x5c7c33144720;  1 drivers
S_0x5c7c32f9b1f0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32f9aff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f9c250_0 .net "in_a", 0 0, L_0x5c7c33145130;  alias, 1 drivers
v0x5c7c32f9c320_0 .net "in_b", 0 0, L_0x5c7c331433b0;  alias, 1 drivers
v0x5c7c32f9c3f0_0 .net "out", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
v0x5c7c32f9c510_0 .net "temp_out", 0 0, L_0x5c7c33144510;  1 drivers
S_0x5c7c32f9b460 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f9b1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144510 .functor NAND 1, L_0x5c7c33145130, L_0x5c7c331433b0, C4<1>, C4<1>;
v0x5c7c32f9b6d0_0 .net "in_a", 0 0, L_0x5c7c33145130;  alias, 1 drivers
v0x5c7c32f9b7b0_0 .net "in_b", 0 0, L_0x5c7c331433b0;  alias, 1 drivers
v0x5c7c32f9b870_0 .net "out", 0 0, L_0x5c7c33144510;  alias, 1 drivers
S_0x5c7c32f9b990 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f9b1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f9c0d0_0 .net "in_a", 0 0, L_0x5c7c33144510;  alias, 1 drivers
v0x5c7c32f9c170_0 .net "out", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
S_0x5c7c32f9bbb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f9b990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331445c0 .functor NAND 1, L_0x5c7c33144510, L_0x5c7c33144510, C4<1>, C4<1>;
v0x5c7c32f9be20_0 .net "in_a", 0 0, L_0x5c7c33144510;  alias, 1 drivers
v0x5c7c32f9bee0_0 .net "in_b", 0 0, L_0x5c7c33144510;  alias, 1 drivers
v0x5c7c32f9bfd0_0 .net "out", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
S_0x5c7c32f9c5d0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32f9aff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f9d5e0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f9d680_0 .net "in_b", 0 0, L_0x5c7c331451d0;  alias, 1 drivers
v0x5c7c32f9d770_0 .net "out", 0 0, L_0x5c7c33144720;  alias, 1 drivers
v0x5c7c32f9d890_0 .net "temp_out", 0 0, L_0x5c7c33144670;  1 drivers
S_0x5c7c32f9c7b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f9c5d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144670 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c331451d0, C4<1>, C4<1>;
v0x5c7c32f9ca20_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f9cae0_0 .net "in_b", 0 0, L_0x5c7c331451d0;  alias, 1 drivers
v0x5c7c32f9cba0_0 .net "out", 0 0, L_0x5c7c33144670;  alias, 1 drivers
S_0x5c7c32f9ccc0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f9c5d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f9d430_0 .net "in_a", 0 0, L_0x5c7c33144670;  alias, 1 drivers
v0x5c7c32f9d4d0_0 .net "out", 0 0, L_0x5c7c33144720;  alias, 1 drivers
S_0x5c7c32f9cee0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f9ccc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144720 .functor NAND 1, L_0x5c7c33144670, L_0x5c7c33144670, C4<1>, C4<1>;
v0x5c7c32f9d150_0 .net "in_a", 0 0, L_0x5c7c33144670;  alias, 1 drivers
v0x5c7c32f9d240_0 .net "in_b", 0 0, L_0x5c7c33144670;  alias, 1 drivers
v0x5c7c32f9d330_0 .net "out", 0 0, L_0x5c7c33144720;  alias, 1 drivers
S_0x5c7c32f9d950 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32f9aff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f9e050_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f9e0f0_0 .net "out", 0 0, L_0x5c7c331433b0;  alias, 1 drivers
S_0x5c7c32f9db20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f9d950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331433b0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32f9dd70_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f9de30_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32f9def0_0 .net "out", 0 0, L_0x5c7c331433b0;  alias, 1 drivers
S_0x5c7c32f9e1f0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32f9aff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fa3ca0_0 .net "branch1_out", 0 0, L_0x5c7c33144930;  1 drivers
v0x5c7c32fa3dd0_0 .net "branch2_out", 0 0, L_0x5c7c33144c50;  1 drivers
v0x5c7c32fa3f20_0 .net "in_a", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
v0x5c7c32fa3ff0_0 .net "in_b", 0 0, L_0x5c7c33144720;  alias, 1 drivers
v0x5c7c32fa4090_0 .net "out", 0 0, L_0x5c7c33144f70;  alias, 1 drivers
v0x5c7c32fa4130_0 .net "temp1_out", 0 0, L_0x5c7c33144880;  1 drivers
v0x5c7c32fa41d0_0 .net "temp2_out", 0 0, L_0x5c7c33144ba0;  1 drivers
v0x5c7c32fa4270_0 .net "temp3_out", 0 0, L_0x5c7c33144ec0;  1 drivers
S_0x5c7c32f9e420 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32f9e1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32f9f4e0_0 .net "in_a", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
v0x5c7c32f9f580_0 .net "in_b", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
v0x5c7c32f9f640_0 .net "out", 0 0, L_0x5c7c33144880;  alias, 1 drivers
v0x5c7c32f9f760_0 .net "temp_out", 0 0, L_0x5c7c331447d0;  1 drivers
S_0x5c7c32f9e690 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f9e420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331447d0 .functor NAND 1, L_0x5c7c331445c0, L_0x5c7c331445c0, C4<1>, C4<1>;
v0x5c7c32f9e900_0 .net "in_a", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
v0x5c7c32f9e9c0_0 .net "in_b", 0 0, L_0x5c7c331445c0;  alias, 1 drivers
v0x5c7c32f9eb10_0 .net "out", 0 0, L_0x5c7c331447d0;  alias, 1 drivers
S_0x5c7c32f9ec10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f9e420;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32f9f330_0 .net "in_a", 0 0, L_0x5c7c331447d0;  alias, 1 drivers
v0x5c7c32f9f3d0_0 .net "out", 0 0, L_0x5c7c33144880;  alias, 1 drivers
S_0x5c7c32f9ede0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32f9ec10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144880 .functor NAND 1, L_0x5c7c331447d0, L_0x5c7c331447d0, C4<1>, C4<1>;
v0x5c7c32f9f050_0 .net "in_a", 0 0, L_0x5c7c331447d0;  alias, 1 drivers
v0x5c7c32f9f140_0 .net "in_b", 0 0, L_0x5c7c331447d0;  alias, 1 drivers
v0x5c7c32f9f230_0 .net "out", 0 0, L_0x5c7c33144880;  alias, 1 drivers
S_0x5c7c32f9f8d0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32f9e1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fa0900_0 .net "in_a", 0 0, L_0x5c7c33144720;  alias, 1 drivers
v0x5c7c32fa09a0_0 .net "in_b", 0 0, L_0x5c7c33144720;  alias, 1 drivers
v0x5c7c32fa0a60_0 .net "out", 0 0, L_0x5c7c33144ba0;  alias, 1 drivers
v0x5c7c32fa0b80_0 .net "temp_out", 0 0, L_0x5c7c33144af0;  1 drivers
S_0x5c7c32f9fab0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32f9f8d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144af0 .functor NAND 1, L_0x5c7c33144720, L_0x5c7c33144720, C4<1>, C4<1>;
v0x5c7c32f9fd20_0 .net "in_a", 0 0, L_0x5c7c33144720;  alias, 1 drivers
v0x5c7c32f9fde0_0 .net "in_b", 0 0, L_0x5c7c33144720;  alias, 1 drivers
v0x5c7c32f9ff30_0 .net "out", 0 0, L_0x5c7c33144af0;  alias, 1 drivers
S_0x5c7c32fa0030 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32f9f8d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa0750_0 .net "in_a", 0 0, L_0x5c7c33144af0;  alias, 1 drivers
v0x5c7c32fa07f0_0 .net "out", 0 0, L_0x5c7c33144ba0;  alias, 1 drivers
S_0x5c7c32fa0200 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa0030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144ba0 .functor NAND 1, L_0x5c7c33144af0, L_0x5c7c33144af0, C4<1>, C4<1>;
v0x5c7c32fa0470_0 .net "in_a", 0 0, L_0x5c7c33144af0;  alias, 1 drivers
v0x5c7c32fa0560_0 .net "in_b", 0 0, L_0x5c7c33144af0;  alias, 1 drivers
v0x5c7c32fa0650_0 .net "out", 0 0, L_0x5c7c33144ba0;  alias, 1 drivers
S_0x5c7c32fa0cf0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32f9e1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fa1d30_0 .net "in_a", 0 0, L_0x5c7c33144930;  alias, 1 drivers
v0x5c7c32fa1e00_0 .net "in_b", 0 0, L_0x5c7c33144c50;  alias, 1 drivers
v0x5c7c32fa1ed0_0 .net "out", 0 0, L_0x5c7c33144ec0;  alias, 1 drivers
v0x5c7c32fa1ff0_0 .net "temp_out", 0 0, L_0x5c7c33144e10;  1 drivers
S_0x5c7c32fa0ed0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fa0cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144e10 .functor NAND 1, L_0x5c7c33144930, L_0x5c7c33144c50, C4<1>, C4<1>;
v0x5c7c32fa1120_0 .net "in_a", 0 0, L_0x5c7c33144930;  alias, 1 drivers
v0x5c7c32fa1200_0 .net "in_b", 0 0, L_0x5c7c33144c50;  alias, 1 drivers
v0x5c7c32fa12c0_0 .net "out", 0 0, L_0x5c7c33144e10;  alias, 1 drivers
S_0x5c7c32fa1410 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fa0cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa1b80_0 .net "in_a", 0 0, L_0x5c7c33144e10;  alias, 1 drivers
v0x5c7c32fa1c20_0 .net "out", 0 0, L_0x5c7c33144ec0;  alias, 1 drivers
S_0x5c7c32fa1630 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa1410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144ec0 .functor NAND 1, L_0x5c7c33144e10, L_0x5c7c33144e10, C4<1>, C4<1>;
v0x5c7c32fa18a0_0 .net "in_a", 0 0, L_0x5c7c33144e10;  alias, 1 drivers
v0x5c7c32fa1990_0 .net "in_b", 0 0, L_0x5c7c33144e10;  alias, 1 drivers
v0x5c7c32fa1a80_0 .net "out", 0 0, L_0x5c7c33144ec0;  alias, 1 drivers
S_0x5c7c32fa2140 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32f9e1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa2870_0 .net "in_a", 0 0, L_0x5c7c33144880;  alias, 1 drivers
v0x5c7c32fa2910_0 .net "out", 0 0, L_0x5c7c33144930;  alias, 1 drivers
S_0x5c7c32fa2310 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa2140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144930 .functor NAND 1, L_0x5c7c33144880, L_0x5c7c33144880, C4<1>, C4<1>;
v0x5c7c32fa2580_0 .net "in_a", 0 0, L_0x5c7c33144880;  alias, 1 drivers
v0x5c7c32fa2640_0 .net "in_b", 0 0, L_0x5c7c33144880;  alias, 1 drivers
v0x5c7c32fa2790_0 .net "out", 0 0, L_0x5c7c33144930;  alias, 1 drivers
S_0x5c7c32fa2a10 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32f9e1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa31e0_0 .net "in_a", 0 0, L_0x5c7c33144ba0;  alias, 1 drivers
v0x5c7c32fa3280_0 .net "out", 0 0, L_0x5c7c33144c50;  alias, 1 drivers
S_0x5c7c32fa2c80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa2a10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144c50 .functor NAND 1, L_0x5c7c33144ba0, L_0x5c7c33144ba0, C4<1>, C4<1>;
v0x5c7c32fa2ef0_0 .net "in_a", 0 0, L_0x5c7c33144ba0;  alias, 1 drivers
v0x5c7c32fa2fb0_0 .net "in_b", 0 0, L_0x5c7c33144ba0;  alias, 1 drivers
v0x5c7c32fa3100_0 .net "out", 0 0, L_0x5c7c33144c50;  alias, 1 drivers
S_0x5c7c32fa3380 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32f9e1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa3b20_0 .net "in_a", 0 0, L_0x5c7c33144ec0;  alias, 1 drivers
v0x5c7c32fa3bc0_0 .net "out", 0 0, L_0x5c7c33144f70;  alias, 1 drivers
S_0x5c7c32fa35a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa3380;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33144f70 .functor NAND 1, L_0x5c7c33144ec0, L_0x5c7c33144ec0, C4<1>, C4<1>;
v0x5c7c32fa3810_0 .net "in_a", 0 0, L_0x5c7c33144ec0;  alias, 1 drivers
v0x5c7c32fa38d0_0 .net "in_b", 0 0, L_0x5c7c33144ec0;  alias, 1 drivers
v0x5c7c32fa3a20_0 .net "out", 0 0, L_0x5c7c33144f70;  alias, 1 drivers
S_0x5c7c32fa4b60 .scope module, "mux_gate8" "Mux" 15 15, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fadec0_0 .net "in_a", 0 0, L_0x5c7c33145fd0;  1 drivers
v0x5c7c32fadf60_0 .net "in_b", 0 0, L_0x5c7c33146070;  1 drivers
v0x5c7c32fae070_0 .net "out", 0 0, L_0x5c7c33145e10;  1 drivers
v0x5c7c32fae110_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fae1b0_0 .net "sel_out", 0 0, L_0x5c7c33145300;  1 drivers
v0x5c7c32fae330_0 .net "temp_a_out", 0 0, L_0x5c7c33145460;  1 drivers
v0x5c7c32fae4e0_0 .net "temp_b_out", 0 0, L_0x5c7c331455c0;  1 drivers
S_0x5c7c32fa4d60 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fa4b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fa5dc0_0 .net "in_a", 0 0, L_0x5c7c33145fd0;  alias, 1 drivers
v0x5c7c32fa5e90_0 .net "in_b", 0 0, L_0x5c7c33145300;  alias, 1 drivers
v0x5c7c32fa5f60_0 .net "out", 0 0, L_0x5c7c33145460;  alias, 1 drivers
v0x5c7c32fa6080_0 .net "temp_out", 0 0, L_0x5c7c331453b0;  1 drivers
S_0x5c7c32fa4fd0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fa4d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331453b0 .functor NAND 1, L_0x5c7c33145fd0, L_0x5c7c33145300, C4<1>, C4<1>;
v0x5c7c32fa5240_0 .net "in_a", 0 0, L_0x5c7c33145fd0;  alias, 1 drivers
v0x5c7c32fa5320_0 .net "in_b", 0 0, L_0x5c7c33145300;  alias, 1 drivers
v0x5c7c32fa53e0_0 .net "out", 0 0, L_0x5c7c331453b0;  alias, 1 drivers
S_0x5c7c32fa5500 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fa4d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa5c40_0 .net "in_a", 0 0, L_0x5c7c331453b0;  alias, 1 drivers
v0x5c7c32fa5ce0_0 .net "out", 0 0, L_0x5c7c33145460;  alias, 1 drivers
S_0x5c7c32fa5720 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa5500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145460 .functor NAND 1, L_0x5c7c331453b0, L_0x5c7c331453b0, C4<1>, C4<1>;
v0x5c7c32fa5990_0 .net "in_a", 0 0, L_0x5c7c331453b0;  alias, 1 drivers
v0x5c7c32fa5a50_0 .net "in_b", 0 0, L_0x5c7c331453b0;  alias, 1 drivers
v0x5c7c32fa5b40_0 .net "out", 0 0, L_0x5c7c33145460;  alias, 1 drivers
S_0x5c7c32fa6140 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fa4b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fa7150_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fa71f0_0 .net "in_b", 0 0, L_0x5c7c33146070;  alias, 1 drivers
v0x5c7c32fa72e0_0 .net "out", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
v0x5c7c32fa7400_0 .net "temp_out", 0 0, L_0x5c7c33145510;  1 drivers
S_0x5c7c32fa6320 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fa6140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145510 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33146070, C4<1>, C4<1>;
v0x5c7c32fa6590_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fa6650_0 .net "in_b", 0 0, L_0x5c7c33146070;  alias, 1 drivers
v0x5c7c32fa6710_0 .net "out", 0 0, L_0x5c7c33145510;  alias, 1 drivers
S_0x5c7c32fa6830 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fa6140;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa6fa0_0 .net "in_a", 0 0, L_0x5c7c33145510;  alias, 1 drivers
v0x5c7c32fa7040_0 .net "out", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
S_0x5c7c32fa6a50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa6830;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331455c0 .functor NAND 1, L_0x5c7c33145510, L_0x5c7c33145510, C4<1>, C4<1>;
v0x5c7c32fa6cc0_0 .net "in_a", 0 0, L_0x5c7c33145510;  alias, 1 drivers
v0x5c7c32fa6db0_0 .net "in_b", 0 0, L_0x5c7c33145510;  alias, 1 drivers
v0x5c7c32fa6ea0_0 .net "out", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
S_0x5c7c32fa74c0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fa4b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa7bc0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fa7c60_0 .net "out", 0 0, L_0x5c7c33145300;  alias, 1 drivers
S_0x5c7c32fa7690 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa74c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145300 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32fa78e0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fa79a0_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fa7a60_0 .net "out", 0 0, L_0x5c7c33145300;  alias, 1 drivers
S_0x5c7c32fa7d60 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fa4b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fad810_0 .net "branch1_out", 0 0, L_0x5c7c331457d0;  1 drivers
v0x5c7c32fad940_0 .net "branch2_out", 0 0, L_0x5c7c33145af0;  1 drivers
v0x5c7c32fada90_0 .net "in_a", 0 0, L_0x5c7c33145460;  alias, 1 drivers
v0x5c7c32fadb60_0 .net "in_b", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
v0x5c7c32fadc00_0 .net "out", 0 0, L_0x5c7c33145e10;  alias, 1 drivers
v0x5c7c32fadca0_0 .net "temp1_out", 0 0, L_0x5c7c33145720;  1 drivers
v0x5c7c32fadd40_0 .net "temp2_out", 0 0, L_0x5c7c33145a40;  1 drivers
v0x5c7c32fadde0_0 .net "temp3_out", 0 0, L_0x5c7c33145d60;  1 drivers
S_0x5c7c32fa7f90 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fa7d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fa9050_0 .net "in_a", 0 0, L_0x5c7c33145460;  alias, 1 drivers
v0x5c7c32fa90f0_0 .net "in_b", 0 0, L_0x5c7c33145460;  alias, 1 drivers
v0x5c7c32fa91b0_0 .net "out", 0 0, L_0x5c7c33145720;  alias, 1 drivers
v0x5c7c32fa92d0_0 .net "temp_out", 0 0, L_0x5c7c33145670;  1 drivers
S_0x5c7c32fa8200 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fa7f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145670 .functor NAND 1, L_0x5c7c33145460, L_0x5c7c33145460, C4<1>, C4<1>;
v0x5c7c32fa8470_0 .net "in_a", 0 0, L_0x5c7c33145460;  alias, 1 drivers
v0x5c7c32fa8530_0 .net "in_b", 0 0, L_0x5c7c33145460;  alias, 1 drivers
v0x5c7c32fa8680_0 .net "out", 0 0, L_0x5c7c33145670;  alias, 1 drivers
S_0x5c7c32fa8780 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fa7f90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fa8ea0_0 .net "in_a", 0 0, L_0x5c7c33145670;  alias, 1 drivers
v0x5c7c32fa8f40_0 .net "out", 0 0, L_0x5c7c33145720;  alias, 1 drivers
S_0x5c7c32fa8950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa8780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145720 .functor NAND 1, L_0x5c7c33145670, L_0x5c7c33145670, C4<1>, C4<1>;
v0x5c7c32fa8bc0_0 .net "in_a", 0 0, L_0x5c7c33145670;  alias, 1 drivers
v0x5c7c32fa8cb0_0 .net "in_b", 0 0, L_0x5c7c33145670;  alias, 1 drivers
v0x5c7c32fa8da0_0 .net "out", 0 0, L_0x5c7c33145720;  alias, 1 drivers
S_0x5c7c32fa9440 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fa7d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32faa470_0 .net "in_a", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
v0x5c7c32faa510_0 .net "in_b", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
v0x5c7c32faa5d0_0 .net "out", 0 0, L_0x5c7c33145a40;  alias, 1 drivers
v0x5c7c32faa6f0_0 .net "temp_out", 0 0, L_0x5c7c33145990;  1 drivers
S_0x5c7c32fa9620 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fa9440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145990 .functor NAND 1, L_0x5c7c331455c0, L_0x5c7c331455c0, C4<1>, C4<1>;
v0x5c7c32fa9890_0 .net "in_a", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
v0x5c7c32fa9950_0 .net "in_b", 0 0, L_0x5c7c331455c0;  alias, 1 drivers
v0x5c7c32fa9aa0_0 .net "out", 0 0, L_0x5c7c33145990;  alias, 1 drivers
S_0x5c7c32fa9ba0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fa9440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32faa2c0_0 .net "in_a", 0 0, L_0x5c7c33145990;  alias, 1 drivers
v0x5c7c32faa360_0 .net "out", 0 0, L_0x5c7c33145a40;  alias, 1 drivers
S_0x5c7c32fa9d70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fa9ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145a40 .functor NAND 1, L_0x5c7c33145990, L_0x5c7c33145990, C4<1>, C4<1>;
v0x5c7c32fa9fe0_0 .net "in_a", 0 0, L_0x5c7c33145990;  alias, 1 drivers
v0x5c7c32faa0d0_0 .net "in_b", 0 0, L_0x5c7c33145990;  alias, 1 drivers
v0x5c7c32faa1c0_0 .net "out", 0 0, L_0x5c7c33145a40;  alias, 1 drivers
S_0x5c7c32faa860 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fa7d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fab8a0_0 .net "in_a", 0 0, L_0x5c7c331457d0;  alias, 1 drivers
v0x5c7c32fab970_0 .net "in_b", 0 0, L_0x5c7c33145af0;  alias, 1 drivers
v0x5c7c32faba40_0 .net "out", 0 0, L_0x5c7c33145d60;  alias, 1 drivers
v0x5c7c32fabb60_0 .net "temp_out", 0 0, L_0x5c7c33145cb0;  1 drivers
S_0x5c7c32faaa40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32faa860;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145cb0 .functor NAND 1, L_0x5c7c331457d0, L_0x5c7c33145af0, C4<1>, C4<1>;
v0x5c7c32faac90_0 .net "in_a", 0 0, L_0x5c7c331457d0;  alias, 1 drivers
v0x5c7c32faad70_0 .net "in_b", 0 0, L_0x5c7c33145af0;  alias, 1 drivers
v0x5c7c32faae30_0 .net "out", 0 0, L_0x5c7c33145cb0;  alias, 1 drivers
S_0x5c7c32faaf80 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32faa860;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fab6f0_0 .net "in_a", 0 0, L_0x5c7c33145cb0;  alias, 1 drivers
v0x5c7c32fab790_0 .net "out", 0 0, L_0x5c7c33145d60;  alias, 1 drivers
S_0x5c7c32fab1a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32faaf80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145d60 .functor NAND 1, L_0x5c7c33145cb0, L_0x5c7c33145cb0, C4<1>, C4<1>;
v0x5c7c32fab410_0 .net "in_a", 0 0, L_0x5c7c33145cb0;  alias, 1 drivers
v0x5c7c32fab500_0 .net "in_b", 0 0, L_0x5c7c33145cb0;  alias, 1 drivers
v0x5c7c32fab5f0_0 .net "out", 0 0, L_0x5c7c33145d60;  alias, 1 drivers
S_0x5c7c32fabcb0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fa7d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fac3e0_0 .net "in_a", 0 0, L_0x5c7c33145720;  alias, 1 drivers
v0x5c7c32fac480_0 .net "out", 0 0, L_0x5c7c331457d0;  alias, 1 drivers
S_0x5c7c32fabe80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fabcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331457d0 .functor NAND 1, L_0x5c7c33145720, L_0x5c7c33145720, C4<1>, C4<1>;
v0x5c7c32fac0f0_0 .net "in_a", 0 0, L_0x5c7c33145720;  alias, 1 drivers
v0x5c7c32fac1b0_0 .net "in_b", 0 0, L_0x5c7c33145720;  alias, 1 drivers
v0x5c7c32fac300_0 .net "out", 0 0, L_0x5c7c331457d0;  alias, 1 drivers
S_0x5c7c32fac580 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fa7d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32facd50_0 .net "in_a", 0 0, L_0x5c7c33145a40;  alias, 1 drivers
v0x5c7c32facdf0_0 .net "out", 0 0, L_0x5c7c33145af0;  alias, 1 drivers
S_0x5c7c32fac7f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fac580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145af0 .functor NAND 1, L_0x5c7c33145a40, L_0x5c7c33145a40, C4<1>, C4<1>;
v0x5c7c32faca60_0 .net "in_a", 0 0, L_0x5c7c33145a40;  alias, 1 drivers
v0x5c7c32facb20_0 .net "in_b", 0 0, L_0x5c7c33145a40;  alias, 1 drivers
v0x5c7c32facc70_0 .net "out", 0 0, L_0x5c7c33145af0;  alias, 1 drivers
S_0x5c7c32facef0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fa7d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fad690_0 .net "in_a", 0 0, L_0x5c7c33145d60;  alias, 1 drivers
v0x5c7c32fad730_0 .net "out", 0 0, L_0x5c7c33145e10;  alias, 1 drivers
S_0x5c7c32fad110 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32facef0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33145e10 .functor NAND 1, L_0x5c7c33145d60, L_0x5c7c33145d60, C4<1>, C4<1>;
v0x5c7c32fad380_0 .net "in_a", 0 0, L_0x5c7c33145d60;  alias, 1 drivers
v0x5c7c32fad440_0 .net "in_b", 0 0, L_0x5c7c33145d60;  alias, 1 drivers
v0x5c7c32fad590_0 .net "out", 0 0, L_0x5c7c33145e10;  alias, 1 drivers
S_0x5c7c32fae6d0 .scope module, "mux_gate9" "Mux" 15 16, 16 3 0, S_0x5c7c32f1b960;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fb7a30_0 .net "in_a", 0 0, L_0x5c7c33146df0;  1 drivers
v0x5c7c32fb7ad0_0 .net "in_b", 0 0, L_0x5c7c33146e90;  1 drivers
v0x5c7c32fb7be0_0 .net "out", 0 0, L_0x5c7c33146c30;  1 drivers
v0x5c7c32fb7c80_0 .net "sel", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fb7d20_0 .net "sel_out", 0 0, L_0x5c7c331461b0;  1 drivers
v0x5c7c32fb7ea0_0 .net "temp_a_out", 0 0, L_0x5c7c33146310;  1 drivers
v0x5c7c32fb8050_0 .net "temp_b_out", 0 0, L_0x5c7c33146470;  1 drivers
S_0x5c7c32fae8d0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fae6d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32faf930_0 .net "in_a", 0 0, L_0x5c7c33146df0;  alias, 1 drivers
v0x5c7c32fafa00_0 .net "in_b", 0 0, L_0x5c7c331461b0;  alias, 1 drivers
v0x5c7c32fafad0_0 .net "out", 0 0, L_0x5c7c33146310;  alias, 1 drivers
v0x5c7c32fafbf0_0 .net "temp_out", 0 0, L_0x5c7c33146260;  1 drivers
S_0x5c7c32faeb40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fae8d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146260 .functor NAND 1, L_0x5c7c33146df0, L_0x5c7c331461b0, C4<1>, C4<1>;
v0x5c7c32faedb0_0 .net "in_a", 0 0, L_0x5c7c33146df0;  alias, 1 drivers
v0x5c7c32faee90_0 .net "in_b", 0 0, L_0x5c7c331461b0;  alias, 1 drivers
v0x5c7c32faef50_0 .net "out", 0 0, L_0x5c7c33146260;  alias, 1 drivers
S_0x5c7c32faf070 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fae8d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32faf7b0_0 .net "in_a", 0 0, L_0x5c7c33146260;  alias, 1 drivers
v0x5c7c32faf850_0 .net "out", 0 0, L_0x5c7c33146310;  alias, 1 drivers
S_0x5c7c32faf290 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32faf070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146310 .functor NAND 1, L_0x5c7c33146260, L_0x5c7c33146260, C4<1>, C4<1>;
v0x5c7c32faf500_0 .net "in_a", 0 0, L_0x5c7c33146260;  alias, 1 drivers
v0x5c7c32faf5c0_0 .net "in_b", 0 0, L_0x5c7c33146260;  alias, 1 drivers
v0x5c7c32faf6b0_0 .net "out", 0 0, L_0x5c7c33146310;  alias, 1 drivers
S_0x5c7c32fafcb0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fae6d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fb0cc0_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fb0d60_0 .net "in_b", 0 0, L_0x5c7c33146e90;  alias, 1 drivers
v0x5c7c32fb0e50_0 .net "out", 0 0, L_0x5c7c33146470;  alias, 1 drivers
v0x5c7c32fb0f70_0 .net "temp_out", 0 0, L_0x5c7c331463c0;  1 drivers
S_0x5c7c32fafe90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fafcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331463c0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c33146e90, C4<1>, C4<1>;
v0x5c7c32fb0100_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fb01c0_0 .net "in_b", 0 0, L_0x5c7c33146e90;  alias, 1 drivers
v0x5c7c32fb0280_0 .net "out", 0 0, L_0x5c7c331463c0;  alias, 1 drivers
S_0x5c7c32fb03a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fafcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb0b10_0 .net "in_a", 0 0, L_0x5c7c331463c0;  alias, 1 drivers
v0x5c7c32fb0bb0_0 .net "out", 0 0, L_0x5c7c33146470;  alias, 1 drivers
S_0x5c7c32fb05c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb03a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146470 .functor NAND 1, L_0x5c7c331463c0, L_0x5c7c331463c0, C4<1>, C4<1>;
v0x5c7c32fb0830_0 .net "in_a", 0 0, L_0x5c7c331463c0;  alias, 1 drivers
v0x5c7c32fb0920_0 .net "in_b", 0 0, L_0x5c7c331463c0;  alias, 1 drivers
v0x5c7c32fb0a10_0 .net "out", 0 0, L_0x5c7c33146470;  alias, 1 drivers
S_0x5c7c32fb1030 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fae6d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb1730_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fb17d0_0 .net "out", 0 0, L_0x5c7c331461b0;  alias, 1 drivers
S_0x5c7c32fb1200 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb1030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331461b0 .functor NAND 1, L_0x5c7c3314c910, L_0x5c7c3314c910, C4<1>, C4<1>;
v0x5c7c32fb1450_0 .net "in_a", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fb1510_0 .net "in_b", 0 0, L_0x5c7c3314c910;  alias, 1 drivers
v0x5c7c32fb15d0_0 .net "out", 0 0, L_0x5c7c331461b0;  alias, 1 drivers
S_0x5c7c32fb18d0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fae6d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fb7380_0 .net "branch1_out", 0 0, L_0x5c7c33146680;  1 drivers
v0x5c7c32fb74b0_0 .net "branch2_out", 0 0, L_0x5c7c331469a0;  1 drivers
v0x5c7c32fb7600_0 .net "in_a", 0 0, L_0x5c7c33146310;  alias, 1 drivers
v0x5c7c32fb76d0_0 .net "in_b", 0 0, L_0x5c7c33146470;  alias, 1 drivers
v0x5c7c32fb7770_0 .net "out", 0 0, L_0x5c7c33146c30;  alias, 1 drivers
v0x5c7c32fb7810_0 .net "temp1_out", 0 0, L_0x5c7c331465d0;  1 drivers
v0x5c7c32fb78b0_0 .net "temp2_out", 0 0, L_0x5c7c331468f0;  1 drivers
v0x5c7c32fb7950_0 .net "temp3_out", 0 0, L_0x5c7c33146b80;  1 drivers
S_0x5c7c32fb1b00 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fb18d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fb2bc0_0 .net "in_a", 0 0, L_0x5c7c33146310;  alias, 1 drivers
v0x5c7c32fb2c60_0 .net "in_b", 0 0, L_0x5c7c33146310;  alias, 1 drivers
v0x5c7c32fb2d20_0 .net "out", 0 0, L_0x5c7c331465d0;  alias, 1 drivers
v0x5c7c32fb2e40_0 .net "temp_out", 0 0, L_0x5c7c33146520;  1 drivers
S_0x5c7c32fb1d70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fb1b00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146520 .functor NAND 1, L_0x5c7c33146310, L_0x5c7c33146310, C4<1>, C4<1>;
v0x5c7c32fb1fe0_0 .net "in_a", 0 0, L_0x5c7c33146310;  alias, 1 drivers
v0x5c7c32fb20a0_0 .net "in_b", 0 0, L_0x5c7c33146310;  alias, 1 drivers
v0x5c7c32fb21f0_0 .net "out", 0 0, L_0x5c7c33146520;  alias, 1 drivers
S_0x5c7c32fb22f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fb1b00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb2a10_0 .net "in_a", 0 0, L_0x5c7c33146520;  alias, 1 drivers
v0x5c7c32fb2ab0_0 .net "out", 0 0, L_0x5c7c331465d0;  alias, 1 drivers
S_0x5c7c32fb24c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb22f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331465d0 .functor NAND 1, L_0x5c7c33146520, L_0x5c7c33146520, C4<1>, C4<1>;
v0x5c7c32fb2730_0 .net "in_a", 0 0, L_0x5c7c33146520;  alias, 1 drivers
v0x5c7c32fb2820_0 .net "in_b", 0 0, L_0x5c7c33146520;  alias, 1 drivers
v0x5c7c32fb2910_0 .net "out", 0 0, L_0x5c7c331465d0;  alias, 1 drivers
S_0x5c7c32fb2fb0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fb18d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fb3fe0_0 .net "in_a", 0 0, L_0x5c7c33146470;  alias, 1 drivers
v0x5c7c32fb4080_0 .net "in_b", 0 0, L_0x5c7c33146470;  alias, 1 drivers
v0x5c7c32fb4140_0 .net "out", 0 0, L_0x5c7c331468f0;  alias, 1 drivers
v0x5c7c32fb4260_0 .net "temp_out", 0 0, L_0x5c7c33146840;  1 drivers
S_0x5c7c32fb3190 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fb2fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146840 .functor NAND 1, L_0x5c7c33146470, L_0x5c7c33146470, C4<1>, C4<1>;
v0x5c7c32fb3400_0 .net "in_a", 0 0, L_0x5c7c33146470;  alias, 1 drivers
v0x5c7c32fb34c0_0 .net "in_b", 0 0, L_0x5c7c33146470;  alias, 1 drivers
v0x5c7c32fb3610_0 .net "out", 0 0, L_0x5c7c33146840;  alias, 1 drivers
S_0x5c7c32fb3710 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fb2fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb3e30_0 .net "in_a", 0 0, L_0x5c7c33146840;  alias, 1 drivers
v0x5c7c32fb3ed0_0 .net "out", 0 0, L_0x5c7c331468f0;  alias, 1 drivers
S_0x5c7c32fb38e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb3710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331468f0 .functor NAND 1, L_0x5c7c33146840, L_0x5c7c33146840, C4<1>, C4<1>;
v0x5c7c32fb3b50_0 .net "in_a", 0 0, L_0x5c7c33146840;  alias, 1 drivers
v0x5c7c32fb3c40_0 .net "in_b", 0 0, L_0x5c7c33146840;  alias, 1 drivers
v0x5c7c32fb3d30_0 .net "out", 0 0, L_0x5c7c331468f0;  alias, 1 drivers
S_0x5c7c32fb43d0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fb18d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fb5410_0 .net "in_a", 0 0, L_0x5c7c33146680;  alias, 1 drivers
v0x5c7c32fb54e0_0 .net "in_b", 0 0, L_0x5c7c331469a0;  alias, 1 drivers
v0x5c7c32fb55b0_0 .net "out", 0 0, L_0x5c7c33146b80;  alias, 1 drivers
v0x5c7c32fb56d0_0 .net "temp_out", 0 0, L_0x5c7c32fb6770;  1 drivers
S_0x5c7c32fb45b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fb43d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c32fb6770 .functor NAND 1, L_0x5c7c33146680, L_0x5c7c331469a0, C4<1>, C4<1>;
v0x5c7c32fb4800_0 .net "in_a", 0 0, L_0x5c7c33146680;  alias, 1 drivers
v0x5c7c32fb48e0_0 .net "in_b", 0 0, L_0x5c7c331469a0;  alias, 1 drivers
v0x5c7c32fb49a0_0 .net "out", 0 0, L_0x5c7c32fb6770;  alias, 1 drivers
S_0x5c7c32fb4af0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fb43d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb5260_0 .net "in_a", 0 0, L_0x5c7c32fb6770;  alias, 1 drivers
v0x5c7c32fb5300_0 .net "out", 0 0, L_0x5c7c33146b80;  alias, 1 drivers
S_0x5c7c32fb4d10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb4af0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146b80 .functor NAND 1, L_0x5c7c32fb6770, L_0x5c7c32fb6770, C4<1>, C4<1>;
v0x5c7c32fb4f80_0 .net "in_a", 0 0, L_0x5c7c32fb6770;  alias, 1 drivers
v0x5c7c32fb5070_0 .net "in_b", 0 0, L_0x5c7c32fb6770;  alias, 1 drivers
v0x5c7c32fb5160_0 .net "out", 0 0, L_0x5c7c33146b80;  alias, 1 drivers
S_0x5c7c32fb5820 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fb18d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb5f50_0 .net "in_a", 0 0, L_0x5c7c331465d0;  alias, 1 drivers
v0x5c7c32fb5ff0_0 .net "out", 0 0, L_0x5c7c33146680;  alias, 1 drivers
S_0x5c7c32fb59f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb5820;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146680 .functor NAND 1, L_0x5c7c331465d0, L_0x5c7c331465d0, C4<1>, C4<1>;
v0x5c7c32fb5c60_0 .net "in_a", 0 0, L_0x5c7c331465d0;  alias, 1 drivers
v0x5c7c32fb5d20_0 .net "in_b", 0 0, L_0x5c7c331465d0;  alias, 1 drivers
v0x5c7c32fb5e70_0 .net "out", 0 0, L_0x5c7c33146680;  alias, 1 drivers
S_0x5c7c32fb60f0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fb18d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb68c0_0 .net "in_a", 0 0, L_0x5c7c331468f0;  alias, 1 drivers
v0x5c7c32fb6960_0 .net "out", 0 0, L_0x5c7c331469a0;  alias, 1 drivers
S_0x5c7c32fb6360 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb60f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331469a0 .functor NAND 1, L_0x5c7c331468f0, L_0x5c7c331468f0, C4<1>, C4<1>;
v0x5c7c32fb65d0_0 .net "in_a", 0 0, L_0x5c7c331468f0;  alias, 1 drivers
v0x5c7c32fb6690_0 .net "in_b", 0 0, L_0x5c7c331468f0;  alias, 1 drivers
v0x5c7c32fb67e0_0 .net "out", 0 0, L_0x5c7c331469a0;  alias, 1 drivers
S_0x5c7c32fb6a60 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fb18d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb7200_0 .net "in_a", 0 0, L_0x5c7c33146b80;  alias, 1 drivers
v0x5c7c32fb72a0_0 .net "out", 0 0, L_0x5c7c33146c30;  alias, 1 drivers
S_0x5c7c32fb6c80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb6a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33146c30 .functor NAND 1, L_0x5c7c33146b80, L_0x5c7c33146b80, C4<1>, C4<1>;
v0x5c7c32fb6ef0_0 .net "in_a", 0 0, L_0x5c7c33146b80;  alias, 1 drivers
v0x5c7c32fb6fb0_0 .net "in_b", 0 0, L_0x5c7c33146b80;  alias, 1 drivers
v0x5c7c32fb7100_0 .net "out", 0 0, L_0x5c7c33146c30;  alias, 1 drivers
S_0x5c7c32fb86e0 .scope module, "mux16_gate2" "Mux16" 14 15, 15 3 0, S_0x5c7c32cac1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "in_a";
    .port_info 1 /INPUT 16 "in_b";
    .port_info 2 /OUTPUT 16 "out";
    .port_info 3 /INPUT 1 "sel";
L_0x5c7c3315b4e0 .functor BUFZ 16, L_0x5c7c3315b440, C4<0000000000000000>, C4<0000000000000000>, C4<0000000000000000>;
v0x5c7c33054950_0 .net "in_a", 15 0, o0x7d2eeb8885c8;  alias, 0 drivers
v0x5c7c33054a50_0 .net "in_b", 15 0, o0x7d2eeb8885f8;  alias, 0 drivers
v0x5c7c33054b30_0 .net "out", 15 0, L_0x5c7c3315b4e0;  alias, 1 drivers
v0x5c7c33054bf0_0 .net "sel", 0 0, L_0x5c7c3315b570;  1 drivers
v0x5c7c33054c90_0 .net/s "tmp_out", 15 0, L_0x5c7c3315b440;  1 drivers
L_0x5c7c3314d680 .part o0x7d2eeb8885c8, 0, 1;
L_0x5c7c3314d740 .part o0x7d2eeb8885f8, 0, 1;
L_0x5c7c3314e4b0 .part o0x7d2eeb8885c8, 1, 1;
L_0x5c7c3314e550 .part o0x7d2eeb8885f8, 1, 1;
L_0x5c7c3314f2a0 .part o0x7d2eeb8885c8, 2, 1;
L_0x5c7c3314f340 .part o0x7d2eeb8885f8, 2, 1;
L_0x5c7c331500f0 .part o0x7d2eeb8885c8, 3, 1;
L_0x5c7c33150190 .part o0x7d2eeb8885f8, 3, 1;
L_0x5c7c33150f00 .part o0x7d2eeb8885c8, 4, 1;
L_0x5c7c33150fa0 .part o0x7d2eeb8885f8, 4, 1;
L_0x5c7c33151d70 .part o0x7d2eeb8885c8, 5, 1;
L_0x5c7c33151e10 .part o0x7d2eeb8885f8, 5, 1;
L_0x5c7c33152bf0 .part o0x7d2eeb8885c8, 6, 1;
L_0x5c7c33152da0 .part o0x7d2eeb8885f8, 6, 1;
L_0x5c7c33153c30 .part o0x7d2eeb8885c8, 7, 1;
L_0x5c7c33153cd0 .part o0x7d2eeb8885f8, 7, 1;
L_0x5c7c33154ad0 .part o0x7d2eeb8885c8, 8, 1;
L_0x5c7c33154b70 .part o0x7d2eeb8885f8, 8, 1;
L_0x5c7c33155980 .part o0x7d2eeb8885c8, 9, 1;
L_0x5c7c33155a20 .part o0x7d2eeb8885f8, 9, 1;
L_0x5c7c33154c10 .part o0x7d2eeb8885c8, 10, 1;
L_0x5c7c33156f80 .part o0x7d2eeb8885f8, 10, 1;
L_0x5c7c33157a30 .part o0x7d2eeb8885c8, 11, 1;
L_0x5c7c33157ad0 .part o0x7d2eeb8885f8, 11, 1;
L_0x5c7c33158590 .part o0x7d2eeb8885c8, 12, 1;
L_0x5c7c33158630 .part o0x7d2eeb8885f8, 12, 1;
L_0x5c7c331591e0 .part o0x7d2eeb8885c8, 13, 1;
L_0x5c7c33159280 .part o0x7d2eeb8885f8, 13, 1;
L_0x5c7c3315a0e0 .part o0x7d2eeb8885c8, 14, 1;
L_0x5c7c3315a390 .part o0x7d2eeb8885f8, 14, 1;
L_0x5c7c3315b1f0 .part o0x7d2eeb8885c8, 15, 1;
L_0x5c7c3315b290 .part o0x7d2eeb8885f8, 15, 1;
LS_0x5c7c3315b440_0_0 .concat8 [ 1 1 1 1], L_0x5c7c3314d4c0, L_0x5c7c3314e2f0, L_0x5c7c3314f0e0, L_0x5c7c3314ff30;
LS_0x5c7c3315b440_0_4 .concat8 [ 1 1 1 1], L_0x5c7c33150d40, L_0x5c7c33151bb0, L_0x5c7c33152a30, L_0x5c7c33153a70;
LS_0x5c7c3315b440_0_8 .concat8 [ 1 1 1 1], L_0x5c7c33154910, L_0x5c7c331557c0, L_0x5c7c33156e00, L_0x5c7c331578b0;
LS_0x5c7c3315b440_0_12 .concat8 [ 1 1 1 1], L_0x5c7c33158410, L_0x5c7c33159020, L_0x5c7c33159f20, L_0x5c7c3315b030;
L_0x5c7c3315b440 .concat8 [ 4 4 4 4], LS_0x5c7c3315b440_0_0, LS_0x5c7c3315b440_0_4, LS_0x5c7c3315b440_0_8, LS_0x5c7c3315b440_0_12;
S_0x5c7c32fb8950 .scope module, "mux_gate0" "Mux" 15 7, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fc1dc0_0 .net "in_a", 0 0, L_0x5c7c3314d680;  1 drivers
v0x5c7c32fc1e60_0 .net "in_b", 0 0, L_0x5c7c3314d740;  1 drivers
v0x5c7c32fc1f70_0 .net "out", 0 0, L_0x5c7c3314d4c0;  1 drivers
v0x5c7c32fc2010_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fc20b0_0 .net "sel_out", 0 0, L_0x5c7c3314c9b0;  1 drivers
v0x5c7c32fc2230_0 .net "temp_a_out", 0 0, L_0x5c7c3314cb10;  1 drivers
v0x5c7c32fc23e0_0 .net "temp_b_out", 0 0, L_0x5c7c3314cc70;  1 drivers
S_0x5c7c32fb8ba0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fb8950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fb9c30_0 .net "in_a", 0 0, L_0x5c7c3314d680;  alias, 1 drivers
v0x5c7c32fb9d00_0 .net "in_b", 0 0, L_0x5c7c3314c9b0;  alias, 1 drivers
v0x5c7c32fb9dd0_0 .net "out", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
v0x5c7c32fb9ef0_0 .net "temp_out", 0 0, L_0x5c7c3314ca60;  1 drivers
S_0x5c7c32fb8e10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fb8ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ca60 .functor NAND 1, L_0x5c7c3314d680, L_0x5c7c3314c9b0, C4<1>, C4<1>;
v0x5c7c32fb9080_0 .net "in_a", 0 0, L_0x5c7c3314d680;  alias, 1 drivers
v0x5c7c32fb9160_0 .net "in_b", 0 0, L_0x5c7c3314c9b0;  alias, 1 drivers
v0x5c7c32fb9220_0 .net "out", 0 0, L_0x5c7c3314ca60;  alias, 1 drivers
S_0x5c7c32fb9340 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fb8ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fb9a80_0 .net "in_a", 0 0, L_0x5c7c3314ca60;  alias, 1 drivers
v0x5c7c32fb9b20_0 .net "out", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
S_0x5c7c32fb9560 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fb9340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314cb10 .functor NAND 1, L_0x5c7c3314ca60, L_0x5c7c3314ca60, C4<1>, C4<1>;
v0x5c7c32fb97d0_0 .net "in_a", 0 0, L_0x5c7c3314ca60;  alias, 1 drivers
v0x5c7c32fb9890_0 .net "in_b", 0 0, L_0x5c7c3314ca60;  alias, 1 drivers
v0x5c7c32fb9980_0 .net "out", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
S_0x5c7c32fb9fb0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fb8950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fbafe0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fbb0b0_0 .net "in_b", 0 0, L_0x5c7c3314d740;  alias, 1 drivers
v0x5c7c32fbb180_0 .net "out", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
v0x5c7c32fbb2a0_0 .net "temp_out", 0 0, L_0x5c7c3314cbc0;  1 drivers
S_0x5c7c32fba190 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fb9fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314cbc0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3314d740, C4<1>, C4<1>;
v0x5c7c32fba400_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fba4e0_0 .net "in_b", 0 0, L_0x5c7c3314d740;  alias, 1 drivers
v0x5c7c32fba5a0_0 .net "out", 0 0, L_0x5c7c3314cbc0;  alias, 1 drivers
S_0x5c7c32fba6c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fb9fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fbae30_0 .net "in_a", 0 0, L_0x5c7c3314cbc0;  alias, 1 drivers
v0x5c7c32fbaed0_0 .net "out", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
S_0x5c7c32fba8e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fba6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314cc70 .functor NAND 1, L_0x5c7c3314cbc0, L_0x5c7c3314cbc0, C4<1>, C4<1>;
v0x5c7c32fbab50_0 .net "in_a", 0 0, L_0x5c7c3314cbc0;  alias, 1 drivers
v0x5c7c32fbac40_0 .net "in_b", 0 0, L_0x5c7c3314cbc0;  alias, 1 drivers
v0x5c7c32fbad30_0 .net "out", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
S_0x5c7c32fbb360 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fb8950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fbba80_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fbbbb0_0 .net "out", 0 0, L_0x5c7c3314c9b0;  alias, 1 drivers
S_0x5c7c32fbb530 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fbb360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314c9b0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fbb780_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fbb890_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fbb950_0 .net "out", 0 0, L_0x5c7c3314c9b0;  alias, 1 drivers
S_0x5c7c32fbbcb0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fb8950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fc1710_0 .net "branch1_out", 0 0, L_0x5c7c3314ce80;  1 drivers
v0x5c7c32fc1840_0 .net "branch2_out", 0 0, L_0x5c7c3314d1a0;  1 drivers
v0x5c7c32fc1990_0 .net "in_a", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
v0x5c7c32fc1a60_0 .net "in_b", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
v0x5c7c32fc1b00_0 .net "out", 0 0, L_0x5c7c3314d4c0;  alias, 1 drivers
v0x5c7c32fc1ba0_0 .net "temp1_out", 0 0, L_0x5c7c3314cdd0;  1 drivers
v0x5c7c32fc1c40_0 .net "temp2_out", 0 0, L_0x5c7c3314d0f0;  1 drivers
v0x5c7c32fc1ce0_0 .net "temp3_out", 0 0, L_0x5c7c3314d410;  1 drivers
S_0x5c7c32fbbe90 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fbbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fbcf50_0 .net "in_a", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
v0x5c7c32fbcff0_0 .net "in_b", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
v0x5c7c32fbd0b0_0 .net "out", 0 0, L_0x5c7c3314cdd0;  alias, 1 drivers
v0x5c7c32fbd1d0_0 .net "temp_out", 0 0, L_0x5c7c3314cd20;  1 drivers
S_0x5c7c32fbc100 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fbbe90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314cd20 .functor NAND 1, L_0x5c7c3314cb10, L_0x5c7c3314cb10, C4<1>, C4<1>;
v0x5c7c32fbc370_0 .net "in_a", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
v0x5c7c32fbc430_0 .net "in_b", 0 0, L_0x5c7c3314cb10;  alias, 1 drivers
v0x5c7c32fbc580_0 .net "out", 0 0, L_0x5c7c3314cd20;  alias, 1 drivers
S_0x5c7c32fbc680 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fbbe90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fbcda0_0 .net "in_a", 0 0, L_0x5c7c3314cd20;  alias, 1 drivers
v0x5c7c32fbce40_0 .net "out", 0 0, L_0x5c7c3314cdd0;  alias, 1 drivers
S_0x5c7c32fbc850 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fbc680;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314cdd0 .functor NAND 1, L_0x5c7c3314cd20, L_0x5c7c3314cd20, C4<1>, C4<1>;
v0x5c7c32fbcac0_0 .net "in_a", 0 0, L_0x5c7c3314cd20;  alias, 1 drivers
v0x5c7c32fbcbb0_0 .net "in_b", 0 0, L_0x5c7c3314cd20;  alias, 1 drivers
v0x5c7c32fbcca0_0 .net "out", 0 0, L_0x5c7c3314cdd0;  alias, 1 drivers
S_0x5c7c32fbd340 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fbbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fbe370_0 .net "in_a", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
v0x5c7c32fbe410_0 .net "in_b", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
v0x5c7c32fbe4d0_0 .net "out", 0 0, L_0x5c7c3314d0f0;  alias, 1 drivers
v0x5c7c32fbe5f0_0 .net "temp_out", 0 0, L_0x5c7c3314d040;  1 drivers
S_0x5c7c32fbd520 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fbd340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d040 .functor NAND 1, L_0x5c7c3314cc70, L_0x5c7c3314cc70, C4<1>, C4<1>;
v0x5c7c32fbd790_0 .net "in_a", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
v0x5c7c32fbd850_0 .net "in_b", 0 0, L_0x5c7c3314cc70;  alias, 1 drivers
v0x5c7c32fbd9a0_0 .net "out", 0 0, L_0x5c7c3314d040;  alias, 1 drivers
S_0x5c7c32fbdaa0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fbd340;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fbe1c0_0 .net "in_a", 0 0, L_0x5c7c3314d040;  alias, 1 drivers
v0x5c7c32fbe260_0 .net "out", 0 0, L_0x5c7c3314d0f0;  alias, 1 drivers
S_0x5c7c32fbdc70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fbdaa0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d0f0 .functor NAND 1, L_0x5c7c3314d040, L_0x5c7c3314d040, C4<1>, C4<1>;
v0x5c7c32fbdee0_0 .net "in_a", 0 0, L_0x5c7c3314d040;  alias, 1 drivers
v0x5c7c32fbdfd0_0 .net "in_b", 0 0, L_0x5c7c3314d040;  alias, 1 drivers
v0x5c7c32fbe0c0_0 .net "out", 0 0, L_0x5c7c3314d0f0;  alias, 1 drivers
S_0x5c7c32fbe760 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fbbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fbf7a0_0 .net "in_a", 0 0, L_0x5c7c3314ce80;  alias, 1 drivers
v0x5c7c32fbf870_0 .net "in_b", 0 0, L_0x5c7c3314d1a0;  alias, 1 drivers
v0x5c7c32fbf940_0 .net "out", 0 0, L_0x5c7c3314d410;  alias, 1 drivers
v0x5c7c32fbfa60_0 .net "temp_out", 0 0, L_0x5c7c3314d360;  1 drivers
S_0x5c7c32fbe940 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fbe760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d360 .functor NAND 1, L_0x5c7c3314ce80, L_0x5c7c3314d1a0, C4<1>, C4<1>;
v0x5c7c32fbeb90_0 .net "in_a", 0 0, L_0x5c7c3314ce80;  alias, 1 drivers
v0x5c7c32fbec70_0 .net "in_b", 0 0, L_0x5c7c3314d1a0;  alias, 1 drivers
v0x5c7c32fbed30_0 .net "out", 0 0, L_0x5c7c3314d360;  alias, 1 drivers
S_0x5c7c32fbee80 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fbe760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fbf5f0_0 .net "in_a", 0 0, L_0x5c7c3314d360;  alias, 1 drivers
v0x5c7c32fbf690_0 .net "out", 0 0, L_0x5c7c3314d410;  alias, 1 drivers
S_0x5c7c32fbf0a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fbee80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d410 .functor NAND 1, L_0x5c7c3314d360, L_0x5c7c3314d360, C4<1>, C4<1>;
v0x5c7c32fbf310_0 .net "in_a", 0 0, L_0x5c7c3314d360;  alias, 1 drivers
v0x5c7c32fbf400_0 .net "in_b", 0 0, L_0x5c7c3314d360;  alias, 1 drivers
v0x5c7c32fbf4f0_0 .net "out", 0 0, L_0x5c7c3314d410;  alias, 1 drivers
S_0x5c7c32fbfbb0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fbbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc02e0_0 .net "in_a", 0 0, L_0x5c7c3314cdd0;  alias, 1 drivers
v0x5c7c32fc0380_0 .net "out", 0 0, L_0x5c7c3314ce80;  alias, 1 drivers
S_0x5c7c32fbfd80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fbfbb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ce80 .functor NAND 1, L_0x5c7c3314cdd0, L_0x5c7c3314cdd0, C4<1>, C4<1>;
v0x5c7c32fbfff0_0 .net "in_a", 0 0, L_0x5c7c3314cdd0;  alias, 1 drivers
v0x5c7c32fc00b0_0 .net "in_b", 0 0, L_0x5c7c3314cdd0;  alias, 1 drivers
v0x5c7c32fc0200_0 .net "out", 0 0, L_0x5c7c3314ce80;  alias, 1 drivers
S_0x5c7c32fc0480 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fbbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc0c50_0 .net "in_a", 0 0, L_0x5c7c3314d0f0;  alias, 1 drivers
v0x5c7c32fc0cf0_0 .net "out", 0 0, L_0x5c7c3314d1a0;  alias, 1 drivers
S_0x5c7c32fc06f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc0480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d1a0 .functor NAND 1, L_0x5c7c3314d0f0, L_0x5c7c3314d0f0, C4<1>, C4<1>;
v0x5c7c32fc0960_0 .net "in_a", 0 0, L_0x5c7c3314d0f0;  alias, 1 drivers
v0x5c7c32fc0a20_0 .net "in_b", 0 0, L_0x5c7c3314d0f0;  alias, 1 drivers
v0x5c7c32fc0b70_0 .net "out", 0 0, L_0x5c7c3314d1a0;  alias, 1 drivers
S_0x5c7c32fc0df0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fbbcb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc1590_0 .net "in_a", 0 0, L_0x5c7c3314d410;  alias, 1 drivers
v0x5c7c32fc1630_0 .net "out", 0 0, L_0x5c7c3314d4c0;  alias, 1 drivers
S_0x5c7c32fc1010 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc0df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d4c0 .functor NAND 1, L_0x5c7c3314d410, L_0x5c7c3314d410, C4<1>, C4<1>;
v0x5c7c32fc1280_0 .net "in_a", 0 0, L_0x5c7c3314d410;  alias, 1 drivers
v0x5c7c32fc1340_0 .net "in_b", 0 0, L_0x5c7c3314d410;  alias, 1 drivers
v0x5c7c32fc1490_0 .net "out", 0 0, L_0x5c7c3314d4c0;  alias, 1 drivers
S_0x5c7c32fc25d0 .scope module, "mux_gate1" "Mux" 15 8, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fcb9b0_0 .net "in_a", 0 0, L_0x5c7c3314e4b0;  1 drivers
v0x5c7c32fcba50_0 .net "in_b", 0 0, L_0x5c7c3314e550;  1 drivers
v0x5c7c32fcbb60_0 .net "out", 0 0, L_0x5c7c3314e2f0;  1 drivers
v0x5c7c32fcbc00_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fcbca0_0 .net "sel_out", 0 0, L_0x5c7c3314d7e0;  1 drivers
v0x5c7c32fcbe20_0 .net "temp_a_out", 0 0, L_0x5c7c3314d940;  1 drivers
v0x5c7c32fcbfd0_0 .net "temp_b_out", 0 0, L_0x5c7c3314daa0;  1 drivers
S_0x5c7c32fc27f0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fc25d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fc3830_0 .net "in_a", 0 0, L_0x5c7c3314e4b0;  alias, 1 drivers
v0x5c7c32fc3900_0 .net "in_b", 0 0, L_0x5c7c3314d7e0;  alias, 1 drivers
v0x5c7c32fc39d0_0 .net "out", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
v0x5c7c32fc3af0_0 .net "temp_out", 0 0, L_0x5c7c3314d890;  1 drivers
S_0x5c7c32fc2a40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fc27f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d890 .functor NAND 1, L_0x5c7c3314e4b0, L_0x5c7c3314d7e0, C4<1>, C4<1>;
v0x5c7c32fc2cb0_0 .net "in_a", 0 0, L_0x5c7c3314e4b0;  alias, 1 drivers
v0x5c7c32fc2d90_0 .net "in_b", 0 0, L_0x5c7c3314d7e0;  alias, 1 drivers
v0x5c7c32fc2e50_0 .net "out", 0 0, L_0x5c7c3314d890;  alias, 1 drivers
S_0x5c7c32fc2f70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fc27f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc36b0_0 .net "in_a", 0 0, L_0x5c7c3314d890;  alias, 1 drivers
v0x5c7c32fc3750_0 .net "out", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
S_0x5c7c32fc3190 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc2f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d940 .functor NAND 1, L_0x5c7c3314d890, L_0x5c7c3314d890, C4<1>, C4<1>;
v0x5c7c32fc3400_0 .net "in_a", 0 0, L_0x5c7c3314d890;  alias, 1 drivers
v0x5c7c32fc34c0_0 .net "in_b", 0 0, L_0x5c7c3314d890;  alias, 1 drivers
v0x5c7c32fc35b0_0 .net "out", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
S_0x5c7c32fc3bb0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fc25d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fc4bc0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fc4c60_0 .net "in_b", 0 0, L_0x5c7c3314e550;  alias, 1 drivers
v0x5c7c32fc4d50_0 .net "out", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
v0x5c7c32fc4e70_0 .net "temp_out", 0 0, L_0x5c7c3314d9f0;  1 drivers
S_0x5c7c32fc3d90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fc3bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d9f0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3314e550, C4<1>, C4<1>;
v0x5c7c32fc4000_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fc40c0_0 .net "in_b", 0 0, L_0x5c7c3314e550;  alias, 1 drivers
v0x5c7c32fc4180_0 .net "out", 0 0, L_0x5c7c3314d9f0;  alias, 1 drivers
S_0x5c7c32fc42a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fc3bb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc4a10_0 .net "in_a", 0 0, L_0x5c7c3314d9f0;  alias, 1 drivers
v0x5c7c32fc4ab0_0 .net "out", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
S_0x5c7c32fc44c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc42a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314daa0 .functor NAND 1, L_0x5c7c3314d9f0, L_0x5c7c3314d9f0, C4<1>, C4<1>;
v0x5c7c32fc4730_0 .net "in_a", 0 0, L_0x5c7c3314d9f0;  alias, 1 drivers
v0x5c7c32fc4820_0 .net "in_b", 0 0, L_0x5c7c3314d9f0;  alias, 1 drivers
v0x5c7c32fc4910_0 .net "out", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
S_0x5c7c32fc4f30 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fc25d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc5740_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fc57e0_0 .net "out", 0 0, L_0x5c7c3314d7e0;  alias, 1 drivers
S_0x5c7c32fc5100 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc4f30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314d7e0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fc5350_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fc5520_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fc55e0_0 .net "out", 0 0, L_0x5c7c3314d7e0;  alias, 1 drivers
S_0x5c7c32fc58e0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fc25d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fcb300_0 .net "branch1_out", 0 0, L_0x5c7c3314dcb0;  1 drivers
v0x5c7c32fcb430_0 .net "branch2_out", 0 0, L_0x5c7c3314dfd0;  1 drivers
v0x5c7c32fcb580_0 .net "in_a", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
v0x5c7c32fcb650_0 .net "in_b", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
v0x5c7c32fcb6f0_0 .net "out", 0 0, L_0x5c7c3314e2f0;  alias, 1 drivers
v0x5c7c32fcb790_0 .net "temp1_out", 0 0, L_0x5c7c3314dc00;  1 drivers
v0x5c7c32fcb830_0 .net "temp2_out", 0 0, L_0x5c7c3314df20;  1 drivers
v0x5c7c32fcb8d0_0 .net "temp3_out", 0 0, L_0x5c7c3314e240;  1 drivers
S_0x5c7c32fc5b10 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fc58e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fc6b40_0 .net "in_a", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
v0x5c7c32fc6be0_0 .net "in_b", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
v0x5c7c32fc6ca0_0 .net "out", 0 0, L_0x5c7c3314dc00;  alias, 1 drivers
v0x5c7c32fc6dc0_0 .net "temp_out", 0 0, L_0x5c7c3314db50;  1 drivers
S_0x5c7c32fc5d80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fc5b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314db50 .functor NAND 1, L_0x5c7c3314d940, L_0x5c7c3314d940, C4<1>, C4<1>;
v0x5c7c32fc5ff0_0 .net "in_a", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
v0x5c7c32fc60b0_0 .net "in_b", 0 0, L_0x5c7c3314d940;  alias, 1 drivers
v0x5c7c32fc6170_0 .net "out", 0 0, L_0x5c7c3314db50;  alias, 1 drivers
S_0x5c7c32fc6270 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fc5b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc6990_0 .net "in_a", 0 0, L_0x5c7c3314db50;  alias, 1 drivers
v0x5c7c32fc6a30_0 .net "out", 0 0, L_0x5c7c3314dc00;  alias, 1 drivers
S_0x5c7c32fc6440 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc6270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314dc00 .functor NAND 1, L_0x5c7c3314db50, L_0x5c7c3314db50, C4<1>, C4<1>;
v0x5c7c32fc66b0_0 .net "in_a", 0 0, L_0x5c7c3314db50;  alias, 1 drivers
v0x5c7c32fc67a0_0 .net "in_b", 0 0, L_0x5c7c3314db50;  alias, 1 drivers
v0x5c7c32fc6890_0 .net "out", 0 0, L_0x5c7c3314dc00;  alias, 1 drivers
S_0x5c7c32fc6f30 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fc58e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fc7f60_0 .net "in_a", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
v0x5c7c32fc8000_0 .net "in_b", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
v0x5c7c32fc80c0_0 .net "out", 0 0, L_0x5c7c3314df20;  alias, 1 drivers
v0x5c7c32fc81e0_0 .net "temp_out", 0 0, L_0x5c7c3314de70;  1 drivers
S_0x5c7c32fc7110 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fc6f30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314de70 .functor NAND 1, L_0x5c7c3314daa0, L_0x5c7c3314daa0, C4<1>, C4<1>;
v0x5c7c32fc7380_0 .net "in_a", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
v0x5c7c32fc7440_0 .net "in_b", 0 0, L_0x5c7c3314daa0;  alias, 1 drivers
v0x5c7c32fc7590_0 .net "out", 0 0, L_0x5c7c3314de70;  alias, 1 drivers
S_0x5c7c32fc7690 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fc6f30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc7db0_0 .net "in_a", 0 0, L_0x5c7c3314de70;  alias, 1 drivers
v0x5c7c32fc7e50_0 .net "out", 0 0, L_0x5c7c3314df20;  alias, 1 drivers
S_0x5c7c32fc7860 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc7690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314df20 .functor NAND 1, L_0x5c7c3314de70, L_0x5c7c3314de70, C4<1>, C4<1>;
v0x5c7c32fc7ad0_0 .net "in_a", 0 0, L_0x5c7c3314de70;  alias, 1 drivers
v0x5c7c32fc7bc0_0 .net "in_b", 0 0, L_0x5c7c3314de70;  alias, 1 drivers
v0x5c7c32fc7cb0_0 .net "out", 0 0, L_0x5c7c3314df20;  alias, 1 drivers
S_0x5c7c32fc8350 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fc58e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fc9390_0 .net "in_a", 0 0, L_0x5c7c3314dcb0;  alias, 1 drivers
v0x5c7c32fc9460_0 .net "in_b", 0 0, L_0x5c7c3314dfd0;  alias, 1 drivers
v0x5c7c32fc9530_0 .net "out", 0 0, L_0x5c7c3314e240;  alias, 1 drivers
v0x5c7c32fc9650_0 .net "temp_out", 0 0, L_0x5c7c3314e190;  1 drivers
S_0x5c7c32fc8530 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fc8350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e190 .functor NAND 1, L_0x5c7c3314dcb0, L_0x5c7c3314dfd0, C4<1>, C4<1>;
v0x5c7c32fc8780_0 .net "in_a", 0 0, L_0x5c7c3314dcb0;  alias, 1 drivers
v0x5c7c32fc8860_0 .net "in_b", 0 0, L_0x5c7c3314dfd0;  alias, 1 drivers
v0x5c7c32fc8920_0 .net "out", 0 0, L_0x5c7c3314e190;  alias, 1 drivers
S_0x5c7c32fc8a70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fc8350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc91e0_0 .net "in_a", 0 0, L_0x5c7c3314e190;  alias, 1 drivers
v0x5c7c32fc9280_0 .net "out", 0 0, L_0x5c7c3314e240;  alias, 1 drivers
S_0x5c7c32fc8c90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc8a70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e240 .functor NAND 1, L_0x5c7c3314e190, L_0x5c7c3314e190, C4<1>, C4<1>;
v0x5c7c32fc8f00_0 .net "in_a", 0 0, L_0x5c7c3314e190;  alias, 1 drivers
v0x5c7c32fc8ff0_0 .net "in_b", 0 0, L_0x5c7c3314e190;  alias, 1 drivers
v0x5c7c32fc90e0_0 .net "out", 0 0, L_0x5c7c3314e240;  alias, 1 drivers
S_0x5c7c32fc97a0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fc58e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fc9ed0_0 .net "in_a", 0 0, L_0x5c7c3314dc00;  alias, 1 drivers
v0x5c7c32fc9f70_0 .net "out", 0 0, L_0x5c7c3314dcb0;  alias, 1 drivers
S_0x5c7c32fc9970 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fc97a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314dcb0 .functor NAND 1, L_0x5c7c3314dc00, L_0x5c7c3314dc00, C4<1>, C4<1>;
v0x5c7c32fc9be0_0 .net "in_a", 0 0, L_0x5c7c3314dc00;  alias, 1 drivers
v0x5c7c32fc9ca0_0 .net "in_b", 0 0, L_0x5c7c3314dc00;  alias, 1 drivers
v0x5c7c32fc9df0_0 .net "out", 0 0, L_0x5c7c3314dcb0;  alias, 1 drivers
S_0x5c7c32fca070 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fc58e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fca840_0 .net "in_a", 0 0, L_0x5c7c3314df20;  alias, 1 drivers
v0x5c7c32fca8e0_0 .net "out", 0 0, L_0x5c7c3314dfd0;  alias, 1 drivers
S_0x5c7c32fca2e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fca070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314dfd0 .functor NAND 1, L_0x5c7c3314df20, L_0x5c7c3314df20, C4<1>, C4<1>;
v0x5c7c32fca550_0 .net "in_a", 0 0, L_0x5c7c3314df20;  alias, 1 drivers
v0x5c7c32fca610_0 .net "in_b", 0 0, L_0x5c7c3314df20;  alias, 1 drivers
v0x5c7c32fca760_0 .net "out", 0 0, L_0x5c7c3314dfd0;  alias, 1 drivers
S_0x5c7c32fca9e0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fc58e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fcb180_0 .net "in_a", 0 0, L_0x5c7c3314e240;  alias, 1 drivers
v0x5c7c32fcb220_0 .net "out", 0 0, L_0x5c7c3314e2f0;  alias, 1 drivers
S_0x5c7c32fcac00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fca9e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e2f0 .functor NAND 1, L_0x5c7c3314e240, L_0x5c7c3314e240, C4<1>, C4<1>;
v0x5c7c32fcae70_0 .net "in_a", 0 0, L_0x5c7c3314e240;  alias, 1 drivers
v0x5c7c32fcaf30_0 .net "in_b", 0 0, L_0x5c7c3314e240;  alias, 1 drivers
v0x5c7c32fcb080_0 .net "out", 0 0, L_0x5c7c3314e2f0;  alias, 1 drivers
S_0x5c7c32fcc1c0 .scope module, "mux_gate10" "Mux" 15 17, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fd5530_0 .net "in_a", 0 0, L_0x5c7c33154c10;  1 drivers
v0x5c7c32fd55d0_0 .net "in_b", 0 0, L_0x5c7c33156f80;  1 drivers
v0x5c7c32fd56e0_0 .net "out", 0 0, L_0x5c7c33156e00;  1 drivers
v0x5c7c32fd5780_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fd5820_0 .net "sel_out", 0 0, L_0x5c7c33155b70;  1 drivers
v0x5c7c32fd59a0_0 .net "temp_a_out", 0 0, L_0x5c7c3301ce50;  1 drivers
v0x5c7c32fd5a40_0 .net "temp_b_out", 0 0, L_0x5c7c3301cfb0;  1 drivers
S_0x5c7c32fcc3c0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fcc1c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fcd430_0 .net "in_a", 0 0, L_0x5c7c33154c10;  alias, 1 drivers
v0x5c7c32fcd500_0 .net "in_b", 0 0, L_0x5c7c33155b70;  alias, 1 drivers
v0x5c7c32fcd5d0_0 .net "out", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
v0x5c7c32fcd6f0_0 .net "temp_out", 0 0, L_0x5c7c3301cda0;  1 drivers
S_0x5c7c32fcc610 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fcc3c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301cda0 .functor NAND 1, L_0x5c7c33154c10, L_0x5c7c33155b70, C4<1>, C4<1>;
v0x5c7c32fcc880_0 .net "in_a", 0 0, L_0x5c7c33154c10;  alias, 1 drivers
v0x5c7c32fcc960_0 .net "in_b", 0 0, L_0x5c7c33155b70;  alias, 1 drivers
v0x5c7c32fcca20_0 .net "out", 0 0, L_0x5c7c3301cda0;  alias, 1 drivers
S_0x5c7c32fccb40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fcc3c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fcd280_0 .net "in_a", 0 0, L_0x5c7c3301cda0;  alias, 1 drivers
v0x5c7c32fcd320_0 .net "out", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
S_0x5c7c32fccd60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fccb40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301ce50 .functor NAND 1, L_0x5c7c3301cda0, L_0x5c7c3301cda0, C4<1>, C4<1>;
v0x5c7c32fccfd0_0 .net "in_a", 0 0, L_0x5c7c3301cda0;  alias, 1 drivers
v0x5c7c32fcd090_0 .net "in_b", 0 0, L_0x5c7c3301cda0;  alias, 1 drivers
v0x5c7c32fcd180_0 .net "out", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
S_0x5c7c32fcd7b0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fcc1c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fce7c0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fce860_0 .net "in_b", 0 0, L_0x5c7c33156f80;  alias, 1 drivers
v0x5c7c32fce950_0 .net "out", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
v0x5c7c32fcea70_0 .net "temp_out", 0 0, L_0x5c7c3301cf00;  1 drivers
S_0x5c7c32fcd990 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fcd7b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301cf00 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33156f80, C4<1>, C4<1>;
v0x5c7c32fcdc00_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fcdcc0_0 .net "in_b", 0 0, L_0x5c7c33156f80;  alias, 1 drivers
v0x5c7c32fcdd80_0 .net "out", 0 0, L_0x5c7c3301cf00;  alias, 1 drivers
S_0x5c7c32fcdea0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fcd7b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fce610_0 .net "in_a", 0 0, L_0x5c7c3301cf00;  alias, 1 drivers
v0x5c7c32fce6b0_0 .net "out", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
S_0x5c7c32fce0c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fcdea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301cfb0 .functor NAND 1, L_0x5c7c3301cf00, L_0x5c7c3301cf00, C4<1>, C4<1>;
v0x5c7c32fce330_0 .net "in_a", 0 0, L_0x5c7c3301cf00;  alias, 1 drivers
v0x5c7c32fce420_0 .net "in_b", 0 0, L_0x5c7c3301cf00;  alias, 1 drivers
v0x5c7c32fce510_0 .net "out", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
S_0x5c7c32fceb30 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fcc1c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fcf230_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fcf2d0_0 .net "out", 0 0, L_0x5c7c33155b70;  alias, 1 drivers
S_0x5c7c32fced00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fceb30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33155b70 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fcef50_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fcf010_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fcf0d0_0 .net "out", 0 0, L_0x5c7c33155b70;  alias, 1 drivers
S_0x5c7c32fcf3d0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fcc1c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fd4e80_0 .net "branch1_out", 0 0, L_0x5c7c3301d1c0;  1 drivers
v0x5c7c32fd4fb0_0 .net "branch2_out", 0 0, L_0x5c7c3301d4e0;  1 drivers
v0x5c7c32fd5100_0 .net "in_a", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
v0x5c7c32fd51d0_0 .net "in_b", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
v0x5c7c32fd5270_0 .net "out", 0 0, L_0x5c7c33156e00;  alias, 1 drivers
v0x5c7c32fd5310_0 .net "temp1_out", 0 0, L_0x5c7c3301d110;  1 drivers
v0x5c7c32fd53b0_0 .net "temp2_out", 0 0, L_0x5c7c3301d430;  1 drivers
v0x5c7c32fd5450_0 .net "temp3_out", 0 0, L_0x5c7c33156d90;  1 drivers
S_0x5c7c32fcf600 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fcf3d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fd06c0_0 .net "in_a", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
v0x5c7c32fd0760_0 .net "in_b", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
v0x5c7c32fd0820_0 .net "out", 0 0, L_0x5c7c3301d110;  alias, 1 drivers
v0x5c7c32fd0940_0 .net "temp_out", 0 0, L_0x5c7c3301d060;  1 drivers
S_0x5c7c32fcf870 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fcf600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301d060 .functor NAND 1, L_0x5c7c3301ce50, L_0x5c7c3301ce50, C4<1>, C4<1>;
v0x5c7c32fcfae0_0 .net "in_a", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
v0x5c7c32fcfba0_0 .net "in_b", 0 0, L_0x5c7c3301ce50;  alias, 1 drivers
v0x5c7c32fcfcf0_0 .net "out", 0 0, L_0x5c7c3301d060;  alias, 1 drivers
S_0x5c7c32fcfdf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fcf600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd0510_0 .net "in_a", 0 0, L_0x5c7c3301d060;  alias, 1 drivers
v0x5c7c32fd05b0_0 .net "out", 0 0, L_0x5c7c3301d110;  alias, 1 drivers
S_0x5c7c32fcffc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fcfdf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301d110 .functor NAND 1, L_0x5c7c3301d060, L_0x5c7c3301d060, C4<1>, C4<1>;
v0x5c7c32fd0230_0 .net "in_a", 0 0, L_0x5c7c3301d060;  alias, 1 drivers
v0x5c7c32fd0320_0 .net "in_b", 0 0, L_0x5c7c3301d060;  alias, 1 drivers
v0x5c7c32fd0410_0 .net "out", 0 0, L_0x5c7c3301d110;  alias, 1 drivers
S_0x5c7c32fd0ab0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fcf3d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fd1ae0_0 .net "in_a", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
v0x5c7c32fd1b80_0 .net "in_b", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
v0x5c7c32fd1c40_0 .net "out", 0 0, L_0x5c7c3301d430;  alias, 1 drivers
v0x5c7c32fd1d60_0 .net "temp_out", 0 0, L_0x5c7c3301d380;  1 drivers
S_0x5c7c32fd0c90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fd0ab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301d380 .functor NAND 1, L_0x5c7c3301cfb0, L_0x5c7c3301cfb0, C4<1>, C4<1>;
v0x5c7c32fd0f00_0 .net "in_a", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
v0x5c7c32fd0fc0_0 .net "in_b", 0 0, L_0x5c7c3301cfb0;  alias, 1 drivers
v0x5c7c32fd1110_0 .net "out", 0 0, L_0x5c7c3301d380;  alias, 1 drivers
S_0x5c7c32fd1210 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fd0ab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd1930_0 .net "in_a", 0 0, L_0x5c7c3301d380;  alias, 1 drivers
v0x5c7c32fd19d0_0 .net "out", 0 0, L_0x5c7c3301d430;  alias, 1 drivers
S_0x5c7c32fd13e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd1210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301d430 .functor NAND 1, L_0x5c7c3301d380, L_0x5c7c3301d380, C4<1>, C4<1>;
v0x5c7c32fd1650_0 .net "in_a", 0 0, L_0x5c7c3301d380;  alias, 1 drivers
v0x5c7c32fd1740_0 .net "in_b", 0 0, L_0x5c7c3301d380;  alias, 1 drivers
v0x5c7c32fd1830_0 .net "out", 0 0, L_0x5c7c3301d430;  alias, 1 drivers
S_0x5c7c32fd1ed0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fcf3d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fd2f10_0 .net "in_a", 0 0, L_0x5c7c3301d1c0;  alias, 1 drivers
v0x5c7c32fd2fe0_0 .net "in_b", 0 0, L_0x5c7c3301d4e0;  alias, 1 drivers
v0x5c7c32fd30b0_0 .net "out", 0 0, L_0x5c7c33156d90;  alias, 1 drivers
v0x5c7c32fd31d0_0 .net "temp_out", 0 0, L_0x5c7c33156d20;  1 drivers
S_0x5c7c32fd20b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fd1ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33156d20 .functor NAND 1, L_0x5c7c3301d1c0, L_0x5c7c3301d4e0, C4<1>, C4<1>;
v0x5c7c32fd2300_0 .net "in_a", 0 0, L_0x5c7c3301d1c0;  alias, 1 drivers
v0x5c7c32fd23e0_0 .net "in_b", 0 0, L_0x5c7c3301d4e0;  alias, 1 drivers
v0x5c7c32fd24a0_0 .net "out", 0 0, L_0x5c7c33156d20;  alias, 1 drivers
S_0x5c7c32fd25f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fd1ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd2d60_0 .net "in_a", 0 0, L_0x5c7c33156d20;  alias, 1 drivers
v0x5c7c32fd2e00_0 .net "out", 0 0, L_0x5c7c33156d90;  alias, 1 drivers
S_0x5c7c32fd2810 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd25f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33156d90 .functor NAND 1, L_0x5c7c33156d20, L_0x5c7c33156d20, C4<1>, C4<1>;
v0x5c7c32fd2a80_0 .net "in_a", 0 0, L_0x5c7c33156d20;  alias, 1 drivers
v0x5c7c32fd2b70_0 .net "in_b", 0 0, L_0x5c7c33156d20;  alias, 1 drivers
v0x5c7c32fd2c60_0 .net "out", 0 0, L_0x5c7c33156d90;  alias, 1 drivers
S_0x5c7c32fd3320 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fcf3d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd3a50_0 .net "in_a", 0 0, L_0x5c7c3301d110;  alias, 1 drivers
v0x5c7c32fd3af0_0 .net "out", 0 0, L_0x5c7c3301d1c0;  alias, 1 drivers
S_0x5c7c32fd34f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd3320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301d1c0 .functor NAND 1, L_0x5c7c3301d110, L_0x5c7c3301d110, C4<1>, C4<1>;
v0x5c7c32fd3760_0 .net "in_a", 0 0, L_0x5c7c3301d110;  alias, 1 drivers
v0x5c7c32fd3820_0 .net "in_b", 0 0, L_0x5c7c3301d110;  alias, 1 drivers
v0x5c7c32fd3970_0 .net "out", 0 0, L_0x5c7c3301d1c0;  alias, 1 drivers
S_0x5c7c32fd3bf0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fcf3d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd43c0_0 .net "in_a", 0 0, L_0x5c7c3301d430;  alias, 1 drivers
v0x5c7c32fd4460_0 .net "out", 0 0, L_0x5c7c3301d4e0;  alias, 1 drivers
S_0x5c7c32fd3e60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd3bf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3301d4e0 .functor NAND 1, L_0x5c7c3301d430, L_0x5c7c3301d430, C4<1>, C4<1>;
v0x5c7c32fd40d0_0 .net "in_a", 0 0, L_0x5c7c3301d430;  alias, 1 drivers
v0x5c7c32fd4190_0 .net "in_b", 0 0, L_0x5c7c3301d430;  alias, 1 drivers
v0x5c7c32fd42e0_0 .net "out", 0 0, L_0x5c7c3301d4e0;  alias, 1 drivers
S_0x5c7c32fd4560 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fcf3d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd4d00_0 .net "in_a", 0 0, L_0x5c7c33156d90;  alias, 1 drivers
v0x5c7c32fd4da0_0 .net "out", 0 0, L_0x5c7c33156e00;  alias, 1 drivers
S_0x5c7c32fd4780 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd4560;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33156e00 .functor NAND 1, L_0x5c7c33156d90, L_0x5c7c33156d90, C4<1>, C4<1>;
v0x5c7c32fd49f0_0 .net "in_a", 0 0, L_0x5c7c33156d90;  alias, 1 drivers
v0x5c7c32fd4ab0_0 .net "in_b", 0 0, L_0x5c7c33156d90;  alias, 1 drivers
v0x5c7c32fd4c00_0 .net "out", 0 0, L_0x5c7c33156e00;  alias, 1 drivers
S_0x5c7c32fd5c30 .scope module, "mux_gate11" "Mux" 15 18, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fdef90_0 .net "in_a", 0 0, L_0x5c7c33157a30;  1 drivers
v0x5c7c32fdf030_0 .net "in_b", 0 0, L_0x5c7c33157ad0;  1 drivers
v0x5c7c32fdf140_0 .net "out", 0 0, L_0x5c7c331578b0;  1 drivers
v0x5c7c32fdf1e0_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fdf280_0 .net "sel_out", 0 0, L_0x5c7c331570e0;  1 drivers
v0x5c7c32fdf400_0 .net "temp_a_out", 0 0, L_0x5c7c331571c0;  1 drivers
v0x5c7c32fdf5b0_0 .net "temp_b_out", 0 0, L_0x5c7c331572a0;  1 drivers
S_0x5c7c32fd5e30 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fd5c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fd6e90_0 .net "in_a", 0 0, L_0x5c7c33157a30;  alias, 1 drivers
v0x5c7c32fd6f60_0 .net "in_b", 0 0, L_0x5c7c331570e0;  alias, 1 drivers
v0x5c7c32fd7030_0 .net "out", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
v0x5c7c32fd7150_0 .net "temp_out", 0 0, L_0x5c7c33157150;  1 drivers
S_0x5c7c32fd60a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fd5e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157150 .functor NAND 1, L_0x5c7c33157a30, L_0x5c7c331570e0, C4<1>, C4<1>;
v0x5c7c32fd6310_0 .net "in_a", 0 0, L_0x5c7c33157a30;  alias, 1 drivers
v0x5c7c32fd63f0_0 .net "in_b", 0 0, L_0x5c7c331570e0;  alias, 1 drivers
v0x5c7c32fd64b0_0 .net "out", 0 0, L_0x5c7c33157150;  alias, 1 drivers
S_0x5c7c32fd65d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fd5e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd6d10_0 .net "in_a", 0 0, L_0x5c7c33157150;  alias, 1 drivers
v0x5c7c32fd6db0_0 .net "out", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
S_0x5c7c32fd67f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd65d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331571c0 .functor NAND 1, L_0x5c7c33157150, L_0x5c7c33157150, C4<1>, C4<1>;
v0x5c7c32fd6a60_0 .net "in_a", 0 0, L_0x5c7c33157150;  alias, 1 drivers
v0x5c7c32fd6b20_0 .net "in_b", 0 0, L_0x5c7c33157150;  alias, 1 drivers
v0x5c7c32fd6c10_0 .net "out", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
S_0x5c7c32fd7210 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fd5c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fd8220_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fd82c0_0 .net "in_b", 0 0, L_0x5c7c33157ad0;  alias, 1 drivers
v0x5c7c32fd83b0_0 .net "out", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
v0x5c7c32fd84d0_0 .net "temp_out", 0 0, L_0x5c7c33157230;  1 drivers
S_0x5c7c32fd73f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fd7210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157230 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33157ad0, C4<1>, C4<1>;
v0x5c7c32fd7660_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fd7720_0 .net "in_b", 0 0, L_0x5c7c33157ad0;  alias, 1 drivers
v0x5c7c32fd77e0_0 .net "out", 0 0, L_0x5c7c33157230;  alias, 1 drivers
S_0x5c7c32fd7900 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fd7210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd8070_0 .net "in_a", 0 0, L_0x5c7c33157230;  alias, 1 drivers
v0x5c7c32fd8110_0 .net "out", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
S_0x5c7c32fd7b20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd7900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331572a0 .functor NAND 1, L_0x5c7c33157230, L_0x5c7c33157230, C4<1>, C4<1>;
v0x5c7c32fd7d90_0 .net "in_a", 0 0, L_0x5c7c33157230;  alias, 1 drivers
v0x5c7c32fd7e80_0 .net "in_b", 0 0, L_0x5c7c33157230;  alias, 1 drivers
v0x5c7c32fd7f70_0 .net "out", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
S_0x5c7c32fd8590 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fd5c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd8c90_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fd8d30_0 .net "out", 0 0, L_0x5c7c331570e0;  alias, 1 drivers
S_0x5c7c32fd8760 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd8590;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331570e0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fd89b0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fd8a70_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fd8b30_0 .net "out", 0 0, L_0x5c7c331570e0;  alias, 1 drivers
S_0x5c7c32fd8e30 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fd5c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fde8e0_0 .net "branch1_out", 0 0, L_0x5c7c331573f0;  1 drivers
v0x5c7c32fdea10_0 .net "branch2_out", 0 0, L_0x5c7c33157650;  1 drivers
v0x5c7c32fdeb60_0 .net "in_a", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
v0x5c7c32fdec30_0 .net "in_b", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
v0x5c7c32fdecd0_0 .net "out", 0 0, L_0x5c7c331578b0;  alias, 1 drivers
v0x5c7c32fded70_0 .net "temp1_out", 0 0, L_0x5c7c33157380;  1 drivers
v0x5c7c32fdee10_0 .net "temp2_out", 0 0, L_0x5c7c331575e0;  1 drivers
v0x5c7c32fdeeb0_0 .net "temp3_out", 0 0, L_0x5c7c33157840;  1 drivers
S_0x5c7c32fd9060 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fd8e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fda120_0 .net "in_a", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
v0x5c7c32fda1c0_0 .net "in_b", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
v0x5c7c32fda280_0 .net "out", 0 0, L_0x5c7c33157380;  alias, 1 drivers
v0x5c7c32fda3a0_0 .net "temp_out", 0 0, L_0x5c7c33157310;  1 drivers
S_0x5c7c32fd92d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fd9060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157310 .functor NAND 1, L_0x5c7c331571c0, L_0x5c7c331571c0, C4<1>, C4<1>;
v0x5c7c32fd9540_0 .net "in_a", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
v0x5c7c32fd9600_0 .net "in_b", 0 0, L_0x5c7c331571c0;  alias, 1 drivers
v0x5c7c32fd9750_0 .net "out", 0 0, L_0x5c7c33157310;  alias, 1 drivers
S_0x5c7c32fd9850 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fd9060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fd9f70_0 .net "in_a", 0 0, L_0x5c7c33157310;  alias, 1 drivers
v0x5c7c32fda010_0 .net "out", 0 0, L_0x5c7c33157380;  alias, 1 drivers
S_0x5c7c32fd9a20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fd9850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157380 .functor NAND 1, L_0x5c7c33157310, L_0x5c7c33157310, C4<1>, C4<1>;
v0x5c7c32fd9c90_0 .net "in_a", 0 0, L_0x5c7c33157310;  alias, 1 drivers
v0x5c7c32fd9d80_0 .net "in_b", 0 0, L_0x5c7c33157310;  alias, 1 drivers
v0x5c7c32fd9e70_0 .net "out", 0 0, L_0x5c7c33157380;  alias, 1 drivers
S_0x5c7c32fda510 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fd8e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fdb540_0 .net "in_a", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
v0x5c7c32fdb5e0_0 .net "in_b", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
v0x5c7c32fdb6a0_0 .net "out", 0 0, L_0x5c7c331575e0;  alias, 1 drivers
v0x5c7c32fdb7c0_0 .net "temp_out", 0 0, L_0x5c7c33157570;  1 drivers
S_0x5c7c32fda6f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fda510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157570 .functor NAND 1, L_0x5c7c331572a0, L_0x5c7c331572a0, C4<1>, C4<1>;
v0x5c7c32fda960_0 .net "in_a", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
v0x5c7c32fdaa20_0 .net "in_b", 0 0, L_0x5c7c331572a0;  alias, 1 drivers
v0x5c7c32fdab70_0 .net "out", 0 0, L_0x5c7c33157570;  alias, 1 drivers
S_0x5c7c32fdac70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fda510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fdb390_0 .net "in_a", 0 0, L_0x5c7c33157570;  alias, 1 drivers
v0x5c7c32fdb430_0 .net "out", 0 0, L_0x5c7c331575e0;  alias, 1 drivers
S_0x5c7c32fdae40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fdac70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331575e0 .functor NAND 1, L_0x5c7c33157570, L_0x5c7c33157570, C4<1>, C4<1>;
v0x5c7c32fdb0b0_0 .net "in_a", 0 0, L_0x5c7c33157570;  alias, 1 drivers
v0x5c7c32fdb1a0_0 .net "in_b", 0 0, L_0x5c7c33157570;  alias, 1 drivers
v0x5c7c32fdb290_0 .net "out", 0 0, L_0x5c7c331575e0;  alias, 1 drivers
S_0x5c7c32fdb930 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fd8e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fdc970_0 .net "in_a", 0 0, L_0x5c7c331573f0;  alias, 1 drivers
v0x5c7c32fdca40_0 .net "in_b", 0 0, L_0x5c7c33157650;  alias, 1 drivers
v0x5c7c32fdcb10_0 .net "out", 0 0, L_0x5c7c33157840;  alias, 1 drivers
v0x5c7c32fdcc30_0 .net "temp_out", 0 0, L_0x5c7c331577d0;  1 drivers
S_0x5c7c32fdbb10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fdb930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331577d0 .functor NAND 1, L_0x5c7c331573f0, L_0x5c7c33157650, C4<1>, C4<1>;
v0x5c7c32fdbd60_0 .net "in_a", 0 0, L_0x5c7c331573f0;  alias, 1 drivers
v0x5c7c32fdbe40_0 .net "in_b", 0 0, L_0x5c7c33157650;  alias, 1 drivers
v0x5c7c32fdbf00_0 .net "out", 0 0, L_0x5c7c331577d0;  alias, 1 drivers
S_0x5c7c32fdc050 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fdb930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fdc7c0_0 .net "in_a", 0 0, L_0x5c7c331577d0;  alias, 1 drivers
v0x5c7c32fdc860_0 .net "out", 0 0, L_0x5c7c33157840;  alias, 1 drivers
S_0x5c7c32fdc270 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fdc050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157840 .functor NAND 1, L_0x5c7c331577d0, L_0x5c7c331577d0, C4<1>, C4<1>;
v0x5c7c32fdc4e0_0 .net "in_a", 0 0, L_0x5c7c331577d0;  alias, 1 drivers
v0x5c7c32fdc5d0_0 .net "in_b", 0 0, L_0x5c7c331577d0;  alias, 1 drivers
v0x5c7c32fdc6c0_0 .net "out", 0 0, L_0x5c7c33157840;  alias, 1 drivers
S_0x5c7c32fdcd80 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fd8e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fdd4b0_0 .net "in_a", 0 0, L_0x5c7c33157380;  alias, 1 drivers
v0x5c7c32fdd550_0 .net "out", 0 0, L_0x5c7c331573f0;  alias, 1 drivers
S_0x5c7c32fdcf50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fdcd80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331573f0 .functor NAND 1, L_0x5c7c33157380, L_0x5c7c33157380, C4<1>, C4<1>;
v0x5c7c32fdd1c0_0 .net "in_a", 0 0, L_0x5c7c33157380;  alias, 1 drivers
v0x5c7c32fdd280_0 .net "in_b", 0 0, L_0x5c7c33157380;  alias, 1 drivers
v0x5c7c32fdd3d0_0 .net "out", 0 0, L_0x5c7c331573f0;  alias, 1 drivers
S_0x5c7c32fdd650 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fd8e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fdde20_0 .net "in_a", 0 0, L_0x5c7c331575e0;  alias, 1 drivers
v0x5c7c32fddec0_0 .net "out", 0 0, L_0x5c7c33157650;  alias, 1 drivers
S_0x5c7c32fdd8c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fdd650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157650 .functor NAND 1, L_0x5c7c331575e0, L_0x5c7c331575e0, C4<1>, C4<1>;
v0x5c7c32fddb30_0 .net "in_a", 0 0, L_0x5c7c331575e0;  alias, 1 drivers
v0x5c7c32fddbf0_0 .net "in_b", 0 0, L_0x5c7c331575e0;  alias, 1 drivers
v0x5c7c32fddd40_0 .net "out", 0 0, L_0x5c7c33157650;  alias, 1 drivers
S_0x5c7c32fddfc0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fd8e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fde760_0 .net "in_a", 0 0, L_0x5c7c33157840;  alias, 1 drivers
v0x5c7c32fde800_0 .net "out", 0 0, L_0x5c7c331578b0;  alias, 1 drivers
S_0x5c7c32fde1e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fddfc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331578b0 .functor NAND 1, L_0x5c7c33157840, L_0x5c7c33157840, C4<1>, C4<1>;
v0x5c7c32fde450_0 .net "in_a", 0 0, L_0x5c7c33157840;  alias, 1 drivers
v0x5c7c32fde510_0 .net "in_b", 0 0, L_0x5c7c33157840;  alias, 1 drivers
v0x5c7c32fde660_0 .net "out", 0 0, L_0x5c7c331578b0;  alias, 1 drivers
S_0x5c7c32fdf7a0 .scope module, "mux_gate12" "Mux" 15 19, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32fe8b20_0 .net "in_a", 0 0, L_0x5c7c33158590;  1 drivers
v0x5c7c32fe8bc0_0 .net "in_b", 0 0, L_0x5c7c33158630;  1 drivers
v0x5c7c32fe8cd0_0 .net "out", 0 0, L_0x5c7c33158410;  1 drivers
v0x5c7c32fe8d70_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fe8e10_0 .net "sel_out", 0 0, L_0x5c7c33157c40;  1 drivers
v0x5c7c32fe8f90_0 .net "temp_a_out", 0 0, L_0x5c7c33157d20;  1 drivers
v0x5c7c32fe9140_0 .net "temp_b_out", 0 0, L_0x5c7c33157e00;  1 drivers
S_0x5c7c32fdf9f0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fdf7a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fe0a50_0 .net "in_a", 0 0, L_0x5c7c33158590;  alias, 1 drivers
v0x5c7c32fe0af0_0 .net "in_b", 0 0, L_0x5c7c33157c40;  alias, 1 drivers
v0x5c7c32fe0bc0_0 .net "out", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
v0x5c7c32fe0ce0_0 .net "temp_out", 0 0, L_0x5c7c33157cb0;  1 drivers
S_0x5c7c32fdfc60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fdf9f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157cb0 .functor NAND 1, L_0x5c7c33158590, L_0x5c7c33157c40, C4<1>, C4<1>;
v0x5c7c32fdfed0_0 .net "in_a", 0 0, L_0x5c7c33158590;  alias, 1 drivers
v0x5c7c32fdffb0_0 .net "in_b", 0 0, L_0x5c7c33157c40;  alias, 1 drivers
v0x5c7c32fe0070_0 .net "out", 0 0, L_0x5c7c33157cb0;  alias, 1 drivers
S_0x5c7c32fe0190 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fdf9f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe08d0_0 .net "in_a", 0 0, L_0x5c7c33157cb0;  alias, 1 drivers
v0x5c7c32fe0970_0 .net "out", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
S_0x5c7c32fe03b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe0190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157d20 .functor NAND 1, L_0x5c7c33157cb0, L_0x5c7c33157cb0, C4<1>, C4<1>;
v0x5c7c32fe0620_0 .net "in_a", 0 0, L_0x5c7c33157cb0;  alias, 1 drivers
v0x5c7c32fe06e0_0 .net "in_b", 0 0, L_0x5c7c33157cb0;  alias, 1 drivers
v0x5c7c32fe07d0_0 .net "out", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
S_0x5c7c32fe0da0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fdf7a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fe1db0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fe1e50_0 .net "in_b", 0 0, L_0x5c7c33158630;  alias, 1 drivers
v0x5c7c32fe1f40_0 .net "out", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
v0x5c7c32fe2060_0 .net "temp_out", 0 0, L_0x5c7c33157d90;  1 drivers
S_0x5c7c32fe0f80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fe0da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157d90 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33158630, C4<1>, C4<1>;
v0x5c7c32fe11f0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fe12b0_0 .net "in_b", 0 0, L_0x5c7c33158630;  alias, 1 drivers
v0x5c7c32fe1370_0 .net "out", 0 0, L_0x5c7c33157d90;  alias, 1 drivers
S_0x5c7c32fe1490 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fe0da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe1c00_0 .net "in_a", 0 0, L_0x5c7c33157d90;  alias, 1 drivers
v0x5c7c32fe1ca0_0 .net "out", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
S_0x5c7c32fe16b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe1490;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157e00 .functor NAND 1, L_0x5c7c33157d90, L_0x5c7c33157d90, C4<1>, C4<1>;
v0x5c7c32fe1920_0 .net "in_a", 0 0, L_0x5c7c33157d90;  alias, 1 drivers
v0x5c7c32fe1a10_0 .net "in_b", 0 0, L_0x5c7c33157d90;  alias, 1 drivers
v0x5c7c32fe1b00_0 .net "out", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
S_0x5c7c32fe2120 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fdf7a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe2820_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fe28c0_0 .net "out", 0 0, L_0x5c7c33157c40;  alias, 1 drivers
S_0x5c7c32fe22f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe2120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157c40 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fe2540_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fe2600_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fe26c0_0 .net "out", 0 0, L_0x5c7c33157c40;  alias, 1 drivers
S_0x5c7c32fe29c0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fdf7a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fe8470_0 .net "branch1_out", 0 0, L_0x5c7c33157f50;  1 drivers
v0x5c7c32fe85a0_0 .net "branch2_out", 0 0, L_0x5c7c331581b0;  1 drivers
v0x5c7c32fe86f0_0 .net "in_a", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
v0x5c7c32fe87c0_0 .net "in_b", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
v0x5c7c32fe8860_0 .net "out", 0 0, L_0x5c7c33158410;  alias, 1 drivers
v0x5c7c32fe8900_0 .net "temp1_out", 0 0, L_0x5c7c33157ee0;  1 drivers
v0x5c7c32fe89a0_0 .net "temp2_out", 0 0, L_0x5c7c33158140;  1 drivers
v0x5c7c32fe8a40_0 .net "temp3_out", 0 0, L_0x5c7c331583a0;  1 drivers
S_0x5c7c32fe2bf0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fe29c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fe3cb0_0 .net "in_a", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
v0x5c7c32fe3d50_0 .net "in_b", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
v0x5c7c32fe3e10_0 .net "out", 0 0, L_0x5c7c33157ee0;  alias, 1 drivers
v0x5c7c32fe3f30_0 .net "temp_out", 0 0, L_0x5c7c33157e70;  1 drivers
S_0x5c7c32fe2e60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fe2bf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157e70 .functor NAND 1, L_0x5c7c33157d20, L_0x5c7c33157d20, C4<1>, C4<1>;
v0x5c7c32fe30d0_0 .net "in_a", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
v0x5c7c32fe3190_0 .net "in_b", 0 0, L_0x5c7c33157d20;  alias, 1 drivers
v0x5c7c32fe32e0_0 .net "out", 0 0, L_0x5c7c33157e70;  alias, 1 drivers
S_0x5c7c32fe33e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fe2bf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe3b00_0 .net "in_a", 0 0, L_0x5c7c33157e70;  alias, 1 drivers
v0x5c7c32fe3ba0_0 .net "out", 0 0, L_0x5c7c33157ee0;  alias, 1 drivers
S_0x5c7c32fe35b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe33e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157ee0 .functor NAND 1, L_0x5c7c33157e70, L_0x5c7c33157e70, C4<1>, C4<1>;
v0x5c7c32fe3820_0 .net "in_a", 0 0, L_0x5c7c33157e70;  alias, 1 drivers
v0x5c7c32fe3910_0 .net "in_b", 0 0, L_0x5c7c33157e70;  alias, 1 drivers
v0x5c7c32fe3a00_0 .net "out", 0 0, L_0x5c7c33157ee0;  alias, 1 drivers
S_0x5c7c32fe40a0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fe29c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fe50d0_0 .net "in_a", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
v0x5c7c32fe5170_0 .net "in_b", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
v0x5c7c32fe5230_0 .net "out", 0 0, L_0x5c7c33158140;  alias, 1 drivers
v0x5c7c32fe5350_0 .net "temp_out", 0 0, L_0x5c7c331580d0;  1 drivers
S_0x5c7c32fe4280 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fe40a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331580d0 .functor NAND 1, L_0x5c7c33157e00, L_0x5c7c33157e00, C4<1>, C4<1>;
v0x5c7c32fe44f0_0 .net "in_a", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
v0x5c7c32fe45b0_0 .net "in_b", 0 0, L_0x5c7c33157e00;  alias, 1 drivers
v0x5c7c32fe4700_0 .net "out", 0 0, L_0x5c7c331580d0;  alias, 1 drivers
S_0x5c7c32fe4800 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fe40a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe4f20_0 .net "in_a", 0 0, L_0x5c7c331580d0;  alias, 1 drivers
v0x5c7c32fe4fc0_0 .net "out", 0 0, L_0x5c7c33158140;  alias, 1 drivers
S_0x5c7c32fe49d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe4800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158140 .functor NAND 1, L_0x5c7c331580d0, L_0x5c7c331580d0, C4<1>, C4<1>;
v0x5c7c32fe4c40_0 .net "in_a", 0 0, L_0x5c7c331580d0;  alias, 1 drivers
v0x5c7c32fe4d30_0 .net "in_b", 0 0, L_0x5c7c331580d0;  alias, 1 drivers
v0x5c7c32fe4e20_0 .net "out", 0 0, L_0x5c7c33158140;  alias, 1 drivers
S_0x5c7c32fe54c0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fe29c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fe6500_0 .net "in_a", 0 0, L_0x5c7c33157f50;  alias, 1 drivers
v0x5c7c32fe65d0_0 .net "in_b", 0 0, L_0x5c7c331581b0;  alias, 1 drivers
v0x5c7c32fe66a0_0 .net "out", 0 0, L_0x5c7c331583a0;  alias, 1 drivers
v0x5c7c32fe67c0_0 .net "temp_out", 0 0, L_0x5c7c33158330;  1 drivers
S_0x5c7c32fe56a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fe54c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158330 .functor NAND 1, L_0x5c7c33157f50, L_0x5c7c331581b0, C4<1>, C4<1>;
v0x5c7c32fe58f0_0 .net "in_a", 0 0, L_0x5c7c33157f50;  alias, 1 drivers
v0x5c7c32fe59d0_0 .net "in_b", 0 0, L_0x5c7c331581b0;  alias, 1 drivers
v0x5c7c32fe5a90_0 .net "out", 0 0, L_0x5c7c33158330;  alias, 1 drivers
S_0x5c7c32fe5be0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fe54c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe6350_0 .net "in_a", 0 0, L_0x5c7c33158330;  alias, 1 drivers
v0x5c7c32fe63f0_0 .net "out", 0 0, L_0x5c7c331583a0;  alias, 1 drivers
S_0x5c7c32fe5e00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe5be0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331583a0 .functor NAND 1, L_0x5c7c33158330, L_0x5c7c33158330, C4<1>, C4<1>;
v0x5c7c32fe6070_0 .net "in_a", 0 0, L_0x5c7c33158330;  alias, 1 drivers
v0x5c7c32fe6160_0 .net "in_b", 0 0, L_0x5c7c33158330;  alias, 1 drivers
v0x5c7c32fe6250_0 .net "out", 0 0, L_0x5c7c331583a0;  alias, 1 drivers
S_0x5c7c32fe6910 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fe29c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe7040_0 .net "in_a", 0 0, L_0x5c7c33157ee0;  alias, 1 drivers
v0x5c7c32fe70e0_0 .net "out", 0 0, L_0x5c7c33157f50;  alias, 1 drivers
S_0x5c7c32fe6ae0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe6910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33157f50 .functor NAND 1, L_0x5c7c33157ee0, L_0x5c7c33157ee0, C4<1>, C4<1>;
v0x5c7c32fe6d50_0 .net "in_a", 0 0, L_0x5c7c33157ee0;  alias, 1 drivers
v0x5c7c32fe6e10_0 .net "in_b", 0 0, L_0x5c7c33157ee0;  alias, 1 drivers
v0x5c7c32fe6f60_0 .net "out", 0 0, L_0x5c7c33157f50;  alias, 1 drivers
S_0x5c7c32fe71e0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fe29c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe79b0_0 .net "in_a", 0 0, L_0x5c7c33158140;  alias, 1 drivers
v0x5c7c32fe7a50_0 .net "out", 0 0, L_0x5c7c331581b0;  alias, 1 drivers
S_0x5c7c32fe7450 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe71e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331581b0 .functor NAND 1, L_0x5c7c33158140, L_0x5c7c33158140, C4<1>, C4<1>;
v0x5c7c32fe76c0_0 .net "in_a", 0 0, L_0x5c7c33158140;  alias, 1 drivers
v0x5c7c32fe7780_0 .net "in_b", 0 0, L_0x5c7c33158140;  alias, 1 drivers
v0x5c7c32fe78d0_0 .net "out", 0 0, L_0x5c7c331581b0;  alias, 1 drivers
S_0x5c7c32fe7b50 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fe29c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fe82f0_0 .net "in_a", 0 0, L_0x5c7c331583a0;  alias, 1 drivers
v0x5c7c32fe8390_0 .net "out", 0 0, L_0x5c7c33158410;  alias, 1 drivers
S_0x5c7c32fe7d70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe7b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158410 .functor NAND 1, L_0x5c7c331583a0, L_0x5c7c331583a0, C4<1>, C4<1>;
v0x5c7c32fe7fe0_0 .net "in_a", 0 0, L_0x5c7c331583a0;  alias, 1 drivers
v0x5c7c32fe80a0_0 .net "in_b", 0 0, L_0x5c7c331583a0;  alias, 1 drivers
v0x5c7c32fe81f0_0 .net "out", 0 0, L_0x5c7c33158410;  alias, 1 drivers
S_0x5c7c32fe9330 .scope module, "mux_gate13" "Mux" 15 20, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32ff2690_0 .net "in_a", 0 0, L_0x5c7c331591e0;  1 drivers
v0x5c7c32ff2730_0 .net "in_b", 0 0, L_0x5c7c33159280;  1 drivers
v0x5c7c32ff2840_0 .net "out", 0 0, L_0x5c7c33159020;  1 drivers
v0x5c7c32ff28e0_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ff2980_0 .net "sel_out", 0 0, L_0x5c7c331587b0;  1 drivers
v0x5c7c32ff2b00_0 .net "temp_a_out", 0 0, L_0x5c7c33158890;  1 drivers
v0x5c7c32ff2cb0_0 .net "temp_b_out", 0 0, L_0x5c7c33158970;  1 drivers
S_0x5c7c32fe9530 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32fe9330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fea590_0 .net "in_a", 0 0, L_0x5c7c331591e0;  alias, 1 drivers
v0x5c7c32fea660_0 .net "in_b", 0 0, L_0x5c7c331587b0;  alias, 1 drivers
v0x5c7c32fea730_0 .net "out", 0 0, L_0x5c7c33158890;  alias, 1 drivers
v0x5c7c32fea850_0 .net "temp_out", 0 0, L_0x5c7c33158820;  1 drivers
S_0x5c7c32fe97a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fe9530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158820 .functor NAND 1, L_0x5c7c331591e0, L_0x5c7c331587b0, C4<1>, C4<1>;
v0x5c7c32fe9a10_0 .net "in_a", 0 0, L_0x5c7c331591e0;  alias, 1 drivers
v0x5c7c32fe9af0_0 .net "in_b", 0 0, L_0x5c7c331587b0;  alias, 1 drivers
v0x5c7c32fe9bb0_0 .net "out", 0 0, L_0x5c7c33158820;  alias, 1 drivers
S_0x5c7c32fe9cd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fe9530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fea410_0 .net "in_a", 0 0, L_0x5c7c33158820;  alias, 1 drivers
v0x5c7c32fea4b0_0 .net "out", 0 0, L_0x5c7c33158890;  alias, 1 drivers
S_0x5c7c32fe9ef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fe9cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158890 .functor NAND 1, L_0x5c7c33158820, L_0x5c7c33158820, C4<1>, C4<1>;
v0x5c7c32fea160_0 .net "in_a", 0 0, L_0x5c7c33158820;  alias, 1 drivers
v0x5c7c32fea220_0 .net "in_b", 0 0, L_0x5c7c33158820;  alias, 1 drivers
v0x5c7c32fea310_0 .net "out", 0 0, L_0x5c7c33158890;  alias, 1 drivers
S_0x5c7c32fea910 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32fe9330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32feb920_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32feb9c0_0 .net "in_b", 0 0, L_0x5c7c33159280;  alias, 1 drivers
v0x5c7c32febab0_0 .net "out", 0 0, L_0x5c7c33158970;  alias, 1 drivers
v0x5c7c32febbd0_0 .net "temp_out", 0 0, L_0x5c7c33158900;  1 drivers
S_0x5c7c32feaaf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fea910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158900 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33159280, C4<1>, C4<1>;
v0x5c7c32fead60_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32feae20_0 .net "in_b", 0 0, L_0x5c7c33159280;  alias, 1 drivers
v0x5c7c32feaee0_0 .net "out", 0 0, L_0x5c7c33158900;  alias, 1 drivers
S_0x5c7c32feb000 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fea910;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32feb770_0 .net "in_a", 0 0, L_0x5c7c33158900;  alias, 1 drivers
v0x5c7c32feb810_0 .net "out", 0 0, L_0x5c7c33158970;  alias, 1 drivers
S_0x5c7c32feb220 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32feb000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158970 .functor NAND 1, L_0x5c7c33158900, L_0x5c7c33158900, C4<1>, C4<1>;
v0x5c7c32feb490_0 .net "in_a", 0 0, L_0x5c7c33158900;  alias, 1 drivers
v0x5c7c32feb580_0 .net "in_b", 0 0, L_0x5c7c33158900;  alias, 1 drivers
v0x5c7c32feb670_0 .net "out", 0 0, L_0x5c7c33158970;  alias, 1 drivers
S_0x5c7c32febc90 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32fe9330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fec390_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fec430_0 .net "out", 0 0, L_0x5c7c331587b0;  alias, 1 drivers
S_0x5c7c32febe60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32febc90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331587b0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fec0b0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fec170_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fec230_0 .net "out", 0 0, L_0x5c7c331587b0;  alias, 1 drivers
S_0x5c7c32fec530 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32fe9330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff1fe0_0 .net "branch1_out", 0 0, L_0x5c7c33158ac0;  1 drivers
v0x5c7c32ff2110_0 .net "branch2_out", 0 0, L_0x5c7c33158d20;  1 drivers
v0x5c7c32ff2260_0 .net "in_a", 0 0, L_0x5c7c33158890;  alias, 1 drivers
v0x5c7c32ff2330_0 .net "in_b", 0 0, L_0x5c7c33158970;  alias, 1 drivers
v0x5c7c32ff23d0_0 .net "out", 0 0, L_0x5c7c33159020;  alias, 1 drivers
v0x5c7c32ff2470_0 .net "temp1_out", 0 0, L_0x5c7c33158a50;  1 drivers
v0x5c7c32ff2510_0 .net "temp2_out", 0 0, L_0x5c7c33158cb0;  1 drivers
v0x5c7c32ff25b0_0 .net "temp3_out", 0 0, L_0x5c7c33158f70;  1 drivers
S_0x5c7c32fec760 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fec530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fed820_0 .net "in_a", 0 0, L_0x5c7c33158890;  alias, 1 drivers
v0x5c7c32fed8c0_0 .net "in_b", 0 0, L_0x5c7c33158890;  alias, 1 drivers
v0x5c7c32fed980_0 .net "out", 0 0, L_0x5c7c33158a50;  alias, 1 drivers
v0x5c7c32fedaa0_0 .net "temp_out", 0 0, L_0x5c7c331589e0;  1 drivers
S_0x5c7c32fec9d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fec760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331589e0 .functor NAND 1, L_0x5c7c33158890, L_0x5c7c33158890, C4<1>, C4<1>;
v0x5c7c32fecc40_0 .net "in_a", 0 0, L_0x5c7c33158890;  alias, 1 drivers
v0x5c7c32fecd00_0 .net "in_b", 0 0, L_0x5c7c33158890;  alias, 1 drivers
v0x5c7c32fece50_0 .net "out", 0 0, L_0x5c7c331589e0;  alias, 1 drivers
S_0x5c7c32fecf50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fec760;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fed670_0 .net "in_a", 0 0, L_0x5c7c331589e0;  alias, 1 drivers
v0x5c7c32fed710_0 .net "out", 0 0, L_0x5c7c33158a50;  alias, 1 drivers
S_0x5c7c32fed120 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fecf50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158a50 .functor NAND 1, L_0x5c7c331589e0, L_0x5c7c331589e0, C4<1>, C4<1>;
v0x5c7c32fed390_0 .net "in_a", 0 0, L_0x5c7c331589e0;  alias, 1 drivers
v0x5c7c32fed480_0 .net "in_b", 0 0, L_0x5c7c331589e0;  alias, 1 drivers
v0x5c7c32fed570_0 .net "out", 0 0, L_0x5c7c33158a50;  alias, 1 drivers
S_0x5c7c32fedc10 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fec530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32feec40_0 .net "in_a", 0 0, L_0x5c7c33158970;  alias, 1 drivers
v0x5c7c32feece0_0 .net "in_b", 0 0, L_0x5c7c33158970;  alias, 1 drivers
v0x5c7c32feeda0_0 .net "out", 0 0, L_0x5c7c33158cb0;  alias, 1 drivers
v0x5c7c32feeec0_0 .net "temp_out", 0 0, L_0x5c7c33158c40;  1 drivers
S_0x5c7c32feddf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fedc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158c40 .functor NAND 1, L_0x5c7c33158970, L_0x5c7c33158970, C4<1>, C4<1>;
v0x5c7c32fee060_0 .net "in_a", 0 0, L_0x5c7c33158970;  alias, 1 drivers
v0x5c7c32fee120_0 .net "in_b", 0 0, L_0x5c7c33158970;  alias, 1 drivers
v0x5c7c32fee270_0 .net "out", 0 0, L_0x5c7c33158c40;  alias, 1 drivers
S_0x5c7c32fee370 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fedc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32feea90_0 .net "in_a", 0 0, L_0x5c7c33158c40;  alias, 1 drivers
v0x5c7c32feeb30_0 .net "out", 0 0, L_0x5c7c33158cb0;  alias, 1 drivers
S_0x5c7c32fee540 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fee370;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158cb0 .functor NAND 1, L_0x5c7c33158c40, L_0x5c7c33158c40, C4<1>, C4<1>;
v0x5c7c32fee7b0_0 .net "in_a", 0 0, L_0x5c7c33158c40;  alias, 1 drivers
v0x5c7c32fee8a0_0 .net "in_b", 0 0, L_0x5c7c33158c40;  alias, 1 drivers
v0x5c7c32fee990_0 .net "out", 0 0, L_0x5c7c33158cb0;  alias, 1 drivers
S_0x5c7c32fef030 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fec530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff0070_0 .net "in_a", 0 0, L_0x5c7c33158ac0;  alias, 1 drivers
v0x5c7c32ff0140_0 .net "in_b", 0 0, L_0x5c7c33158d20;  alias, 1 drivers
v0x5c7c32ff0210_0 .net "out", 0 0, L_0x5c7c33158f70;  alias, 1 drivers
v0x5c7c32ff0330_0 .net "temp_out", 0 0, L_0x5c7c33158ec0;  1 drivers
S_0x5c7c32fef210 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fef030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158ec0 .functor NAND 1, L_0x5c7c33158ac0, L_0x5c7c33158d20, C4<1>, C4<1>;
v0x5c7c32fef460_0 .net "in_a", 0 0, L_0x5c7c33158ac0;  alias, 1 drivers
v0x5c7c32fef540_0 .net "in_b", 0 0, L_0x5c7c33158d20;  alias, 1 drivers
v0x5c7c32fef600_0 .net "out", 0 0, L_0x5c7c33158ec0;  alias, 1 drivers
S_0x5c7c32fef750 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fef030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fefec0_0 .net "in_a", 0 0, L_0x5c7c33158ec0;  alias, 1 drivers
v0x5c7c32feff60_0 .net "out", 0 0, L_0x5c7c33158f70;  alias, 1 drivers
S_0x5c7c32fef970 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fef750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158f70 .functor NAND 1, L_0x5c7c33158ec0, L_0x5c7c33158ec0, C4<1>, C4<1>;
v0x5c7c32fefbe0_0 .net "in_a", 0 0, L_0x5c7c33158ec0;  alias, 1 drivers
v0x5c7c32fefcd0_0 .net "in_b", 0 0, L_0x5c7c33158ec0;  alias, 1 drivers
v0x5c7c32fefdc0_0 .net "out", 0 0, L_0x5c7c33158f70;  alias, 1 drivers
S_0x5c7c32ff0480 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fec530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff0bb0_0 .net "in_a", 0 0, L_0x5c7c33158a50;  alias, 1 drivers
v0x5c7c32ff0c50_0 .net "out", 0 0, L_0x5c7c33158ac0;  alias, 1 drivers
S_0x5c7c32ff0650 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff0480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158ac0 .functor NAND 1, L_0x5c7c33158a50, L_0x5c7c33158a50, C4<1>, C4<1>;
v0x5c7c32ff08c0_0 .net "in_a", 0 0, L_0x5c7c33158a50;  alias, 1 drivers
v0x5c7c32ff0980_0 .net "in_b", 0 0, L_0x5c7c33158a50;  alias, 1 drivers
v0x5c7c32ff0ad0_0 .net "out", 0 0, L_0x5c7c33158ac0;  alias, 1 drivers
S_0x5c7c32ff0d50 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fec530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff1520_0 .net "in_a", 0 0, L_0x5c7c33158cb0;  alias, 1 drivers
v0x5c7c32ff15c0_0 .net "out", 0 0, L_0x5c7c33158d20;  alias, 1 drivers
S_0x5c7c32ff0fc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff0d50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33158d20 .functor NAND 1, L_0x5c7c33158cb0, L_0x5c7c33158cb0, C4<1>, C4<1>;
v0x5c7c32ff1230_0 .net "in_a", 0 0, L_0x5c7c33158cb0;  alias, 1 drivers
v0x5c7c32ff12f0_0 .net "in_b", 0 0, L_0x5c7c33158cb0;  alias, 1 drivers
v0x5c7c32ff1440_0 .net "out", 0 0, L_0x5c7c33158d20;  alias, 1 drivers
S_0x5c7c32ff16c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fec530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff1e60_0 .net "in_a", 0 0, L_0x5c7c33158f70;  alias, 1 drivers
v0x5c7c32ff1f00_0 .net "out", 0 0, L_0x5c7c33159020;  alias, 1 drivers
S_0x5c7c32ff18e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff16c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159020 .functor NAND 1, L_0x5c7c33158f70, L_0x5c7c33158f70, C4<1>, C4<1>;
v0x5c7c32ff1b50_0 .net "in_a", 0 0, L_0x5c7c33158f70;  alias, 1 drivers
v0x5c7c32ff1c10_0 .net "in_b", 0 0, L_0x5c7c33158f70;  alias, 1 drivers
v0x5c7c32ff1d60_0 .net "out", 0 0, L_0x5c7c33159020;  alias, 1 drivers
S_0x5c7c32ff2ea0 .scope module, "mux_gate14" "Mux" 15 21, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c32ffc200_0 .net "in_a", 0 0, L_0x5c7c3315a0e0;  1 drivers
v0x5c7c32ffc2a0_0 .net "in_b", 0 0, L_0x5c7c3315a390;  1 drivers
v0x5c7c32ffc3b0_0 .net "out", 0 0, L_0x5c7c33159f20;  1 drivers
v0x5c7c32ffc450_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ffc4f0_0 .net "sel_out", 0 0, L_0x5c7c33159410;  1 drivers
v0x5c7c32ffc670_0 .net "temp_a_out", 0 0, L_0x5c7c33159570;  1 drivers
v0x5c7c32ffc820_0 .net "temp_b_out", 0 0, L_0x5c7c331596d0;  1 drivers
S_0x5c7c32ff30a0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32ff2ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff4100_0 .net "in_a", 0 0, L_0x5c7c3315a0e0;  alias, 1 drivers
v0x5c7c32ff41d0_0 .net "in_b", 0 0, L_0x5c7c33159410;  alias, 1 drivers
v0x5c7c32ff42a0_0 .net "out", 0 0, L_0x5c7c33159570;  alias, 1 drivers
v0x5c7c32ff43c0_0 .net "temp_out", 0 0, L_0x5c7c331594c0;  1 drivers
S_0x5c7c32ff3310 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ff30a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331594c0 .functor NAND 1, L_0x5c7c3315a0e0, L_0x5c7c33159410, C4<1>, C4<1>;
v0x5c7c32ff3580_0 .net "in_a", 0 0, L_0x5c7c3315a0e0;  alias, 1 drivers
v0x5c7c32ff3660_0 .net "in_b", 0 0, L_0x5c7c33159410;  alias, 1 drivers
v0x5c7c32ff3720_0 .net "out", 0 0, L_0x5c7c331594c0;  alias, 1 drivers
S_0x5c7c32ff3840 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ff30a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff3f80_0 .net "in_a", 0 0, L_0x5c7c331594c0;  alias, 1 drivers
v0x5c7c32ff4020_0 .net "out", 0 0, L_0x5c7c33159570;  alias, 1 drivers
S_0x5c7c32ff3a60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff3840;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159570 .functor NAND 1, L_0x5c7c331594c0, L_0x5c7c331594c0, C4<1>, C4<1>;
v0x5c7c32ff3cd0_0 .net "in_a", 0 0, L_0x5c7c331594c0;  alias, 1 drivers
v0x5c7c32ff3d90_0 .net "in_b", 0 0, L_0x5c7c331594c0;  alias, 1 drivers
v0x5c7c32ff3e80_0 .net "out", 0 0, L_0x5c7c33159570;  alias, 1 drivers
S_0x5c7c32ff4480 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32ff2ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff5490_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ff5530_0 .net "in_b", 0 0, L_0x5c7c3315a390;  alias, 1 drivers
v0x5c7c32ff5620_0 .net "out", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
v0x5c7c32ff5740_0 .net "temp_out", 0 0, L_0x5c7c33159620;  1 drivers
S_0x5c7c32ff4660 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ff4480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159620 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315a390, C4<1>, C4<1>;
v0x5c7c32ff48d0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ff4990_0 .net "in_b", 0 0, L_0x5c7c3315a390;  alias, 1 drivers
v0x5c7c32ff4a50_0 .net "out", 0 0, L_0x5c7c33159620;  alias, 1 drivers
S_0x5c7c32ff4b70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ff4480;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff52e0_0 .net "in_a", 0 0, L_0x5c7c33159620;  alias, 1 drivers
v0x5c7c32ff5380_0 .net "out", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
S_0x5c7c32ff4d90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff4b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331596d0 .functor NAND 1, L_0x5c7c33159620, L_0x5c7c33159620, C4<1>, C4<1>;
v0x5c7c32ff5000_0 .net "in_a", 0 0, L_0x5c7c33159620;  alias, 1 drivers
v0x5c7c32ff50f0_0 .net "in_b", 0 0, L_0x5c7c33159620;  alias, 1 drivers
v0x5c7c32ff51e0_0 .net "out", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
S_0x5c7c32ff5800 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32ff2ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff5f00_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ff5fa0_0 .net "out", 0 0, L_0x5c7c33159410;  alias, 1 drivers
S_0x5c7c32ff59d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff5800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159410 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32ff5c20_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ff5ce0_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ff5da0_0 .net "out", 0 0, L_0x5c7c33159410;  alias, 1 drivers
S_0x5c7c32ff60a0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32ff2ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ffbb50_0 .net "branch1_out", 0 0, L_0x5c7c331598e0;  1 drivers
v0x5c7c32ffbc80_0 .net "branch2_out", 0 0, L_0x5c7c33159c00;  1 drivers
v0x5c7c32ffbdd0_0 .net "in_a", 0 0, L_0x5c7c33159570;  alias, 1 drivers
v0x5c7c32ffbea0_0 .net "in_b", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
v0x5c7c32ffbf40_0 .net "out", 0 0, L_0x5c7c33159f20;  alias, 1 drivers
v0x5c7c32ffbfe0_0 .net "temp1_out", 0 0, L_0x5c7c33159830;  1 drivers
v0x5c7c32ffc080_0 .net "temp2_out", 0 0, L_0x5c7c33159b50;  1 drivers
v0x5c7c32ffc120_0 .net "temp3_out", 0 0, L_0x5c7c33159e70;  1 drivers
S_0x5c7c32ff62d0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32ff60a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff7390_0 .net "in_a", 0 0, L_0x5c7c33159570;  alias, 1 drivers
v0x5c7c32ff7430_0 .net "in_b", 0 0, L_0x5c7c33159570;  alias, 1 drivers
v0x5c7c32ff74f0_0 .net "out", 0 0, L_0x5c7c33159830;  alias, 1 drivers
v0x5c7c32ff7610_0 .net "temp_out", 0 0, L_0x5c7c33159780;  1 drivers
S_0x5c7c32ff6540 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ff62d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159780 .functor NAND 1, L_0x5c7c33159570, L_0x5c7c33159570, C4<1>, C4<1>;
v0x5c7c32ff67b0_0 .net "in_a", 0 0, L_0x5c7c33159570;  alias, 1 drivers
v0x5c7c32ff6870_0 .net "in_b", 0 0, L_0x5c7c33159570;  alias, 1 drivers
v0x5c7c32ff69c0_0 .net "out", 0 0, L_0x5c7c33159780;  alias, 1 drivers
S_0x5c7c32ff6ac0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ff62d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff71e0_0 .net "in_a", 0 0, L_0x5c7c33159780;  alias, 1 drivers
v0x5c7c32ff7280_0 .net "out", 0 0, L_0x5c7c33159830;  alias, 1 drivers
S_0x5c7c32ff6c90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff6ac0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159830 .functor NAND 1, L_0x5c7c33159780, L_0x5c7c33159780, C4<1>, C4<1>;
v0x5c7c32ff6f00_0 .net "in_a", 0 0, L_0x5c7c33159780;  alias, 1 drivers
v0x5c7c32ff6ff0_0 .net "in_b", 0 0, L_0x5c7c33159780;  alias, 1 drivers
v0x5c7c32ff70e0_0 .net "out", 0 0, L_0x5c7c33159830;  alias, 1 drivers
S_0x5c7c32ff7780 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32ff60a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff87b0_0 .net "in_a", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
v0x5c7c32ff8850_0 .net "in_b", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
v0x5c7c32ff8910_0 .net "out", 0 0, L_0x5c7c33159b50;  alias, 1 drivers
v0x5c7c32ff8a30_0 .net "temp_out", 0 0, L_0x5c7c33159aa0;  1 drivers
S_0x5c7c32ff7960 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ff7780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159aa0 .functor NAND 1, L_0x5c7c331596d0, L_0x5c7c331596d0, C4<1>, C4<1>;
v0x5c7c32ff7bd0_0 .net "in_a", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
v0x5c7c32ff7c90_0 .net "in_b", 0 0, L_0x5c7c331596d0;  alias, 1 drivers
v0x5c7c32ff7de0_0 .net "out", 0 0, L_0x5c7c33159aa0;  alias, 1 drivers
S_0x5c7c32ff7ee0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ff7780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff8600_0 .net "in_a", 0 0, L_0x5c7c33159aa0;  alias, 1 drivers
v0x5c7c32ff86a0_0 .net "out", 0 0, L_0x5c7c33159b50;  alias, 1 drivers
S_0x5c7c32ff80b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff7ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159b50 .functor NAND 1, L_0x5c7c33159aa0, L_0x5c7c33159aa0, C4<1>, C4<1>;
v0x5c7c32ff8320_0 .net "in_a", 0 0, L_0x5c7c33159aa0;  alias, 1 drivers
v0x5c7c32ff8410_0 .net "in_b", 0 0, L_0x5c7c33159aa0;  alias, 1 drivers
v0x5c7c32ff8500_0 .net "out", 0 0, L_0x5c7c33159b50;  alias, 1 drivers
S_0x5c7c32ff8ba0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32ff60a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ff9be0_0 .net "in_a", 0 0, L_0x5c7c331598e0;  alias, 1 drivers
v0x5c7c32ff9cb0_0 .net "in_b", 0 0, L_0x5c7c33159c00;  alias, 1 drivers
v0x5c7c32ff9d80_0 .net "out", 0 0, L_0x5c7c33159e70;  alias, 1 drivers
v0x5c7c32ff9ea0_0 .net "temp_out", 0 0, L_0x5c7c33159dc0;  1 drivers
S_0x5c7c32ff8d80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ff8ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159dc0 .functor NAND 1, L_0x5c7c331598e0, L_0x5c7c33159c00, C4<1>, C4<1>;
v0x5c7c32ff8fd0_0 .net "in_a", 0 0, L_0x5c7c331598e0;  alias, 1 drivers
v0x5c7c32ff90b0_0 .net "in_b", 0 0, L_0x5c7c33159c00;  alias, 1 drivers
v0x5c7c32ff9170_0 .net "out", 0 0, L_0x5c7c33159dc0;  alias, 1 drivers
S_0x5c7c32ff92c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ff8ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ff9a30_0 .net "in_a", 0 0, L_0x5c7c33159dc0;  alias, 1 drivers
v0x5c7c32ff9ad0_0 .net "out", 0 0, L_0x5c7c33159e70;  alias, 1 drivers
S_0x5c7c32ff94e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff92c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159e70 .functor NAND 1, L_0x5c7c33159dc0, L_0x5c7c33159dc0, C4<1>, C4<1>;
v0x5c7c32ff9750_0 .net "in_a", 0 0, L_0x5c7c33159dc0;  alias, 1 drivers
v0x5c7c32ff9840_0 .net "in_b", 0 0, L_0x5c7c33159dc0;  alias, 1 drivers
v0x5c7c32ff9930_0 .net "out", 0 0, L_0x5c7c33159e70;  alias, 1 drivers
S_0x5c7c32ff9ff0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32ff60a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ffa720_0 .net "in_a", 0 0, L_0x5c7c33159830;  alias, 1 drivers
v0x5c7c32ffa7c0_0 .net "out", 0 0, L_0x5c7c331598e0;  alias, 1 drivers
S_0x5c7c32ffa1c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ff9ff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331598e0 .functor NAND 1, L_0x5c7c33159830, L_0x5c7c33159830, C4<1>, C4<1>;
v0x5c7c32ffa430_0 .net "in_a", 0 0, L_0x5c7c33159830;  alias, 1 drivers
v0x5c7c32ffa4f0_0 .net "in_b", 0 0, L_0x5c7c33159830;  alias, 1 drivers
v0x5c7c32ffa640_0 .net "out", 0 0, L_0x5c7c331598e0;  alias, 1 drivers
S_0x5c7c32ffa8c0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32ff60a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ffb090_0 .net "in_a", 0 0, L_0x5c7c33159b50;  alias, 1 drivers
v0x5c7c32ffb130_0 .net "out", 0 0, L_0x5c7c33159c00;  alias, 1 drivers
S_0x5c7c32ffab30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ffa8c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159c00 .functor NAND 1, L_0x5c7c33159b50, L_0x5c7c33159b50, C4<1>, C4<1>;
v0x5c7c32ffada0_0 .net "in_a", 0 0, L_0x5c7c33159b50;  alias, 1 drivers
v0x5c7c32ffae60_0 .net "in_b", 0 0, L_0x5c7c33159b50;  alias, 1 drivers
v0x5c7c32ffafb0_0 .net "out", 0 0, L_0x5c7c33159c00;  alias, 1 drivers
S_0x5c7c32ffb230 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32ff60a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ffb9d0_0 .net "in_a", 0 0, L_0x5c7c33159e70;  alias, 1 drivers
v0x5c7c32ffba70_0 .net "out", 0 0, L_0x5c7c33159f20;  alias, 1 drivers
S_0x5c7c32ffb450 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ffb230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33159f20 .functor NAND 1, L_0x5c7c33159e70, L_0x5c7c33159e70, C4<1>, C4<1>;
v0x5c7c32ffb6c0_0 .net "in_a", 0 0, L_0x5c7c33159e70;  alias, 1 drivers
v0x5c7c32ffb780_0 .net "in_b", 0 0, L_0x5c7c33159e70;  alias, 1 drivers
v0x5c7c32ffb8d0_0 .net "out", 0 0, L_0x5c7c33159f20;  alias, 1 drivers
S_0x5c7c32ffca10 .scope module, "mux_gate15" "Mux" 15 22, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33005d70_0 .net "in_a", 0 0, L_0x5c7c3315b1f0;  1 drivers
v0x5c7c33005e10_0 .net "in_b", 0 0, L_0x5c7c3315b290;  1 drivers
v0x5c7c33005f20_0 .net "out", 0 0, L_0x5c7c3315b030;  1 drivers
v0x5c7c33005fc0_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33006060_0 .net "sel_out", 0 0, L_0x5c7c3315a740;  1 drivers
v0x5c7c330061e0_0 .net "temp_a_out", 0 0, L_0x5c7c3315a8a0;  1 drivers
v0x5c7c33006390_0 .net "temp_b_out", 0 0, L_0x5c7c3315aa00;  1 drivers
S_0x5c7c32ffcc10 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c32ffca10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32ffdc70_0 .net "in_a", 0 0, L_0x5c7c3315b1f0;  alias, 1 drivers
v0x5c7c32ffdd40_0 .net "in_b", 0 0, L_0x5c7c3315a740;  alias, 1 drivers
v0x5c7c32ffde10_0 .net "out", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
v0x5c7c32ffdf30_0 .net "temp_out", 0 0, L_0x5c7c3315a7f0;  1 drivers
S_0x5c7c32ffce80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ffcc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315a7f0 .functor NAND 1, L_0x5c7c3315b1f0, L_0x5c7c3315a740, C4<1>, C4<1>;
v0x5c7c32ffd0f0_0 .net "in_a", 0 0, L_0x5c7c3315b1f0;  alias, 1 drivers
v0x5c7c32ffd1d0_0 .net "in_b", 0 0, L_0x5c7c3315a740;  alias, 1 drivers
v0x5c7c32ffd290_0 .net "out", 0 0, L_0x5c7c3315a7f0;  alias, 1 drivers
S_0x5c7c32ffd3b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ffcc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ffdaf0_0 .net "in_a", 0 0, L_0x5c7c3315a7f0;  alias, 1 drivers
v0x5c7c32ffdb90_0 .net "out", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
S_0x5c7c32ffd5d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ffd3b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315a8a0 .functor NAND 1, L_0x5c7c3315a7f0, L_0x5c7c3315a7f0, C4<1>, C4<1>;
v0x5c7c32ffd840_0 .net "in_a", 0 0, L_0x5c7c3315a7f0;  alias, 1 drivers
v0x5c7c32ffd900_0 .net "in_b", 0 0, L_0x5c7c3315a7f0;  alias, 1 drivers
v0x5c7c32ffd9f0_0 .net "out", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
S_0x5c7c32ffdff0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c32ffca10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c32fff000_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fff0a0_0 .net "in_b", 0 0, L_0x5c7c3315b290;  alias, 1 drivers
v0x5c7c32fff190_0 .net "out", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
v0x5c7c32fff2b0_0 .net "temp_out", 0 0, L_0x5c7c3315a950;  1 drivers
S_0x5c7c32ffe1d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32ffdff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315a950 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b290, C4<1>, C4<1>;
v0x5c7c32ffe440_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32ffe500_0 .net "in_b", 0 0, L_0x5c7c3315b290;  alias, 1 drivers
v0x5c7c32ffe5c0_0 .net "out", 0 0, L_0x5c7c3315a950;  alias, 1 drivers
S_0x5c7c32ffe6e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32ffdff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32ffee50_0 .net "in_a", 0 0, L_0x5c7c3315a950;  alias, 1 drivers
v0x5c7c32ffeef0_0 .net "out", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
S_0x5c7c32ffe900 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32ffe6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315aa00 .functor NAND 1, L_0x5c7c3315a950, L_0x5c7c3315a950, C4<1>, C4<1>;
v0x5c7c32ffeb70_0 .net "in_a", 0 0, L_0x5c7c3315a950;  alias, 1 drivers
v0x5c7c32ffec60_0 .net "in_b", 0 0, L_0x5c7c3315a950;  alias, 1 drivers
v0x5c7c32ffed50_0 .net "out", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
S_0x5c7c32fff370 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c32ffca10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c32fffa70_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fffb10_0 .net "out", 0 0, L_0x5c7c3315a740;  alias, 1 drivers
S_0x5c7c32fff540 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c32fff370;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315a740 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c32fff790_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fff850_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c32fff910_0 .net "out", 0 0, L_0x5c7c3315a740;  alias, 1 drivers
S_0x5c7c32fffc10 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c32ffca10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330056c0_0 .net "branch1_out", 0 0, L_0x5c7c3315ac10;  1 drivers
v0x5c7c330057f0_0 .net "branch2_out", 0 0, L_0x5c7c3315ae20;  1 drivers
v0x5c7c33005940_0 .net "in_a", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
v0x5c7c33005a10_0 .net "in_b", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
v0x5c7c33005ab0_0 .net "out", 0 0, L_0x5c7c3315b030;  alias, 1 drivers
v0x5c7c33005b50_0 .net "temp1_out", 0 0, L_0x5c7c3315ab60;  1 drivers
v0x5c7c33005bf0_0 .net "temp2_out", 0 0, L_0x5c7c3315ad70;  1 drivers
v0x5c7c33005c90_0 .net "temp3_out", 0 0, L_0x5c7c3315af80;  1 drivers
S_0x5c7c32fffe40 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c32fffc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33000f00_0 .net "in_a", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
v0x5c7c33000fa0_0 .net "in_b", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
v0x5c7c33001060_0 .net "out", 0 0, L_0x5c7c3315ab60;  alias, 1 drivers
v0x5c7c33001180_0 .net "temp_out", 0 0, L_0x5c7c3315aab0;  1 drivers
S_0x5c7c330000b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c32fffe40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315aab0 .functor NAND 1, L_0x5c7c3315a8a0, L_0x5c7c3315a8a0, C4<1>, C4<1>;
v0x5c7c33000320_0 .net "in_a", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
v0x5c7c330003e0_0 .net "in_b", 0 0, L_0x5c7c3315a8a0;  alias, 1 drivers
v0x5c7c33000530_0 .net "out", 0 0, L_0x5c7c3315aab0;  alias, 1 drivers
S_0x5c7c33000630 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c32fffe40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33000d50_0 .net "in_a", 0 0, L_0x5c7c3315aab0;  alias, 1 drivers
v0x5c7c33000df0_0 .net "out", 0 0, L_0x5c7c3315ab60;  alias, 1 drivers
S_0x5c7c33000800 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33000630;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ab60 .functor NAND 1, L_0x5c7c3315aab0, L_0x5c7c3315aab0, C4<1>, C4<1>;
v0x5c7c33000a70_0 .net "in_a", 0 0, L_0x5c7c3315aab0;  alias, 1 drivers
v0x5c7c33000b60_0 .net "in_b", 0 0, L_0x5c7c3315aab0;  alias, 1 drivers
v0x5c7c33000c50_0 .net "out", 0 0, L_0x5c7c3315ab60;  alias, 1 drivers
S_0x5c7c330012f0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c32fffc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33002320_0 .net "in_a", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
v0x5c7c330023c0_0 .net "in_b", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
v0x5c7c33002480_0 .net "out", 0 0, L_0x5c7c3315ad70;  alias, 1 drivers
v0x5c7c330025a0_0 .net "temp_out", 0 0, L_0x5c7c3315acc0;  1 drivers
S_0x5c7c330014d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330012f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315acc0 .functor NAND 1, L_0x5c7c3315aa00, L_0x5c7c3315aa00, C4<1>, C4<1>;
v0x5c7c33001740_0 .net "in_a", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
v0x5c7c33001800_0 .net "in_b", 0 0, L_0x5c7c3315aa00;  alias, 1 drivers
v0x5c7c33001950_0 .net "out", 0 0, L_0x5c7c3315acc0;  alias, 1 drivers
S_0x5c7c33001a50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330012f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33002170_0 .net "in_a", 0 0, L_0x5c7c3315acc0;  alias, 1 drivers
v0x5c7c33002210_0 .net "out", 0 0, L_0x5c7c3315ad70;  alias, 1 drivers
S_0x5c7c33001c20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33001a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ad70 .functor NAND 1, L_0x5c7c3315acc0, L_0x5c7c3315acc0, C4<1>, C4<1>;
v0x5c7c33001e90_0 .net "in_a", 0 0, L_0x5c7c3315acc0;  alias, 1 drivers
v0x5c7c33001f80_0 .net "in_b", 0 0, L_0x5c7c3315acc0;  alias, 1 drivers
v0x5c7c33002070_0 .net "out", 0 0, L_0x5c7c3315ad70;  alias, 1 drivers
S_0x5c7c33002710 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c32fffc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33003750_0 .net "in_a", 0 0, L_0x5c7c3315ac10;  alias, 1 drivers
v0x5c7c33003820_0 .net "in_b", 0 0, L_0x5c7c3315ae20;  alias, 1 drivers
v0x5c7c330038f0_0 .net "out", 0 0, L_0x5c7c3315af80;  alias, 1 drivers
v0x5c7c33003a10_0 .net "temp_out", 0 0, L_0x5c7c3315aed0;  1 drivers
S_0x5c7c330028f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33002710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315aed0 .functor NAND 1, L_0x5c7c3315ac10, L_0x5c7c3315ae20, C4<1>, C4<1>;
v0x5c7c33002b40_0 .net "in_a", 0 0, L_0x5c7c3315ac10;  alias, 1 drivers
v0x5c7c33002c20_0 .net "in_b", 0 0, L_0x5c7c3315ae20;  alias, 1 drivers
v0x5c7c33002ce0_0 .net "out", 0 0, L_0x5c7c3315aed0;  alias, 1 drivers
S_0x5c7c33002e30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33002710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330035a0_0 .net "in_a", 0 0, L_0x5c7c3315aed0;  alias, 1 drivers
v0x5c7c33003640_0 .net "out", 0 0, L_0x5c7c3315af80;  alias, 1 drivers
S_0x5c7c33003050 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33002e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315af80 .functor NAND 1, L_0x5c7c3315aed0, L_0x5c7c3315aed0, C4<1>, C4<1>;
v0x5c7c330032c0_0 .net "in_a", 0 0, L_0x5c7c3315aed0;  alias, 1 drivers
v0x5c7c330033b0_0 .net "in_b", 0 0, L_0x5c7c3315aed0;  alias, 1 drivers
v0x5c7c330034a0_0 .net "out", 0 0, L_0x5c7c3315af80;  alias, 1 drivers
S_0x5c7c33003b60 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c32fffc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33004290_0 .net "in_a", 0 0, L_0x5c7c3315ab60;  alias, 1 drivers
v0x5c7c33004330_0 .net "out", 0 0, L_0x5c7c3315ac10;  alias, 1 drivers
S_0x5c7c33003d30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33003b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ac10 .functor NAND 1, L_0x5c7c3315ab60, L_0x5c7c3315ab60, C4<1>, C4<1>;
v0x5c7c33003fa0_0 .net "in_a", 0 0, L_0x5c7c3315ab60;  alias, 1 drivers
v0x5c7c33004060_0 .net "in_b", 0 0, L_0x5c7c3315ab60;  alias, 1 drivers
v0x5c7c330041b0_0 .net "out", 0 0, L_0x5c7c3315ac10;  alias, 1 drivers
S_0x5c7c33004430 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c32fffc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33004c00_0 .net "in_a", 0 0, L_0x5c7c3315ad70;  alias, 1 drivers
v0x5c7c33004ca0_0 .net "out", 0 0, L_0x5c7c3315ae20;  alias, 1 drivers
S_0x5c7c330046a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33004430;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ae20 .functor NAND 1, L_0x5c7c3315ad70, L_0x5c7c3315ad70, C4<1>, C4<1>;
v0x5c7c33004910_0 .net "in_a", 0 0, L_0x5c7c3315ad70;  alias, 1 drivers
v0x5c7c330049d0_0 .net "in_b", 0 0, L_0x5c7c3315ad70;  alias, 1 drivers
v0x5c7c33004b20_0 .net "out", 0 0, L_0x5c7c3315ae20;  alias, 1 drivers
S_0x5c7c33004da0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c32fffc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33005540_0 .net "in_a", 0 0, L_0x5c7c3315af80;  alias, 1 drivers
v0x5c7c330055e0_0 .net "out", 0 0, L_0x5c7c3315b030;  alias, 1 drivers
S_0x5c7c33004fc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33004da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b030 .functor NAND 1, L_0x5c7c3315af80, L_0x5c7c3315af80, C4<1>, C4<1>;
v0x5c7c33005230_0 .net "in_a", 0 0, L_0x5c7c3315af80;  alias, 1 drivers
v0x5c7c330052f0_0 .net "in_b", 0 0, L_0x5c7c3315af80;  alias, 1 drivers
v0x5c7c33005440_0 .net "out", 0 0, L_0x5c7c3315b030;  alias, 1 drivers
S_0x5c7c33006580 .scope module, "mux_gate2" "Mux" 15 9, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c3300f920_0 .net "in_a", 0 0, L_0x5c7c3314f2a0;  1 drivers
v0x5c7c3300f9c0_0 .net "in_b", 0 0, L_0x5c7c3314f340;  1 drivers
v0x5c7c3300fad0_0 .net "out", 0 0, L_0x5c7c3314f0e0;  1 drivers
v0x5c7c3300fb70_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3300fc10_0 .net "sel_out", 0 0, L_0x5c7c3314e5f0;  1 drivers
v0x5c7c3300fd90_0 .net "temp_a_out", 0 0, L_0x5c7c3314e730;  1 drivers
v0x5c7c3300ff40_0 .net "temp_b_out", 0 0, L_0x5c7c3314e890;  1 drivers
S_0x5c7c33006780 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33006580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33007790_0 .net "in_a", 0 0, L_0x5c7c3314f2a0;  alias, 1 drivers
v0x5c7c33007860_0 .net "in_b", 0 0, L_0x5c7c3314e5f0;  alias, 1 drivers
v0x5c7c33007930_0 .net "out", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
v0x5c7c33007a50_0 .net "temp_out", 0 0, L_0x5c7c3314e680;  1 drivers
S_0x5c7c330069a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33006780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e680 .functor NAND 1, L_0x5c7c3314f2a0, L_0x5c7c3314e5f0, C4<1>, C4<1>;
v0x5c7c33006c10_0 .net "in_a", 0 0, L_0x5c7c3314f2a0;  alias, 1 drivers
v0x5c7c33006cf0_0 .net "in_b", 0 0, L_0x5c7c3314e5f0;  alias, 1 drivers
v0x5c7c33006db0_0 .net "out", 0 0, L_0x5c7c3314e680;  alias, 1 drivers
S_0x5c7c33006ed0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33006780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33007610_0 .net "in_a", 0 0, L_0x5c7c3314e680;  alias, 1 drivers
v0x5c7c330076b0_0 .net "out", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
S_0x5c7c330070f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33006ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e730 .functor NAND 1, L_0x5c7c3314e680, L_0x5c7c3314e680, C4<1>, C4<1>;
v0x5c7c33007360_0 .net "in_a", 0 0, L_0x5c7c3314e680;  alias, 1 drivers
v0x5c7c33007420_0 .net "in_b", 0 0, L_0x5c7c3314e680;  alias, 1 drivers
v0x5c7c33007510_0 .net "out", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
S_0x5c7c33007b10 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33006580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33008b20_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33008bc0_0 .net "in_b", 0 0, L_0x5c7c3314f340;  alias, 1 drivers
v0x5c7c33008cb0_0 .net "out", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
v0x5c7c33008dd0_0 .net "temp_out", 0 0, L_0x5c7c3314e7e0;  1 drivers
S_0x5c7c33007cf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33007b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e7e0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3314f340, C4<1>, C4<1>;
v0x5c7c33007f60_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33008020_0 .net "in_b", 0 0, L_0x5c7c3314f340;  alias, 1 drivers
v0x5c7c330080e0_0 .net "out", 0 0, L_0x5c7c3314e7e0;  alias, 1 drivers
S_0x5c7c33008200 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33007b10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33008970_0 .net "in_a", 0 0, L_0x5c7c3314e7e0;  alias, 1 drivers
v0x5c7c33008a10_0 .net "out", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
S_0x5c7c33008420 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33008200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e890 .functor NAND 1, L_0x5c7c3314e7e0, L_0x5c7c3314e7e0, C4<1>, C4<1>;
v0x5c7c33008690_0 .net "in_a", 0 0, L_0x5c7c3314e7e0;  alias, 1 drivers
v0x5c7c33008780_0 .net "in_b", 0 0, L_0x5c7c3314e7e0;  alias, 1 drivers
v0x5c7c33008870_0 .net "out", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
S_0x5c7c33008f20 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33006580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33009620_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330096c0_0 .net "out", 0 0, L_0x5c7c3314e5f0;  alias, 1 drivers
S_0x5c7c330090f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33008f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e5f0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c33009340_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33009400_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330094c0_0 .net "out", 0 0, L_0x5c7c3314e5f0;  alias, 1 drivers
S_0x5c7c330097c0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33006580;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3300f270_0 .net "branch1_out", 0 0, L_0x5c7c3314eaa0;  1 drivers
v0x5c7c3300f3a0_0 .net "branch2_out", 0 0, L_0x5c7c3314edc0;  1 drivers
v0x5c7c3300f4f0_0 .net "in_a", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
v0x5c7c3300f5c0_0 .net "in_b", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
v0x5c7c3300f660_0 .net "out", 0 0, L_0x5c7c3314f0e0;  alias, 1 drivers
v0x5c7c3300f700_0 .net "temp1_out", 0 0, L_0x5c7c3314e9f0;  1 drivers
v0x5c7c3300f7a0_0 .net "temp2_out", 0 0, L_0x5c7c3314ed10;  1 drivers
v0x5c7c3300f840_0 .net "temp3_out", 0 0, L_0x5c7c3314f030;  1 drivers
S_0x5c7c330099f0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330097c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3300aab0_0 .net "in_a", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
v0x5c7c3300ab50_0 .net "in_b", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
v0x5c7c3300ac10_0 .net "out", 0 0, L_0x5c7c3314e9f0;  alias, 1 drivers
v0x5c7c3300ad30_0 .net "temp_out", 0 0, L_0x5c7c3314e940;  1 drivers
S_0x5c7c33009c60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330099f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e940 .functor NAND 1, L_0x5c7c3314e730, L_0x5c7c3314e730, C4<1>, C4<1>;
v0x5c7c33009ed0_0 .net "in_a", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
v0x5c7c33009f90_0 .net "in_b", 0 0, L_0x5c7c3314e730;  alias, 1 drivers
v0x5c7c3300a0e0_0 .net "out", 0 0, L_0x5c7c3314e940;  alias, 1 drivers
S_0x5c7c3300a1e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330099f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3300a900_0 .net "in_a", 0 0, L_0x5c7c3314e940;  alias, 1 drivers
v0x5c7c3300a9a0_0 .net "out", 0 0, L_0x5c7c3314e9f0;  alias, 1 drivers
S_0x5c7c3300a3b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3300a1e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314e9f0 .functor NAND 1, L_0x5c7c3314e940, L_0x5c7c3314e940, C4<1>, C4<1>;
v0x5c7c3300a620_0 .net "in_a", 0 0, L_0x5c7c3314e940;  alias, 1 drivers
v0x5c7c3300a710_0 .net "in_b", 0 0, L_0x5c7c3314e940;  alias, 1 drivers
v0x5c7c3300a800_0 .net "out", 0 0, L_0x5c7c3314e9f0;  alias, 1 drivers
S_0x5c7c3300aea0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330097c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3300bed0_0 .net "in_a", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
v0x5c7c3300bf70_0 .net "in_b", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
v0x5c7c3300c030_0 .net "out", 0 0, L_0x5c7c3314ed10;  alias, 1 drivers
v0x5c7c3300c150_0 .net "temp_out", 0 0, L_0x5c7c3314ec60;  1 drivers
S_0x5c7c3300b080 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3300aea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ec60 .functor NAND 1, L_0x5c7c3314e890, L_0x5c7c3314e890, C4<1>, C4<1>;
v0x5c7c3300b2f0_0 .net "in_a", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
v0x5c7c3300b3b0_0 .net "in_b", 0 0, L_0x5c7c3314e890;  alias, 1 drivers
v0x5c7c3300b500_0 .net "out", 0 0, L_0x5c7c3314ec60;  alias, 1 drivers
S_0x5c7c3300b600 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3300aea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3300bd20_0 .net "in_a", 0 0, L_0x5c7c3314ec60;  alias, 1 drivers
v0x5c7c3300bdc0_0 .net "out", 0 0, L_0x5c7c3314ed10;  alias, 1 drivers
S_0x5c7c3300b7d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3300b600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ed10 .functor NAND 1, L_0x5c7c3314ec60, L_0x5c7c3314ec60, C4<1>, C4<1>;
v0x5c7c3300ba40_0 .net "in_a", 0 0, L_0x5c7c3314ec60;  alias, 1 drivers
v0x5c7c3300bb30_0 .net "in_b", 0 0, L_0x5c7c3314ec60;  alias, 1 drivers
v0x5c7c3300bc20_0 .net "out", 0 0, L_0x5c7c3314ed10;  alias, 1 drivers
S_0x5c7c3300c2c0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330097c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3300d300_0 .net "in_a", 0 0, L_0x5c7c3314eaa0;  alias, 1 drivers
v0x5c7c3300d3d0_0 .net "in_b", 0 0, L_0x5c7c3314edc0;  alias, 1 drivers
v0x5c7c3300d4a0_0 .net "out", 0 0, L_0x5c7c3314f030;  alias, 1 drivers
v0x5c7c3300d5c0_0 .net "temp_out", 0 0, L_0x5c7c3314ef80;  1 drivers
S_0x5c7c3300c4a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3300c2c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ef80 .functor NAND 1, L_0x5c7c3314eaa0, L_0x5c7c3314edc0, C4<1>, C4<1>;
v0x5c7c3300c6f0_0 .net "in_a", 0 0, L_0x5c7c3314eaa0;  alias, 1 drivers
v0x5c7c3300c7d0_0 .net "in_b", 0 0, L_0x5c7c3314edc0;  alias, 1 drivers
v0x5c7c3300c890_0 .net "out", 0 0, L_0x5c7c3314ef80;  alias, 1 drivers
S_0x5c7c3300c9e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3300c2c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3300d150_0 .net "in_a", 0 0, L_0x5c7c3314ef80;  alias, 1 drivers
v0x5c7c3300d1f0_0 .net "out", 0 0, L_0x5c7c3314f030;  alias, 1 drivers
S_0x5c7c3300cc00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3300c9e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f030 .functor NAND 1, L_0x5c7c3314ef80, L_0x5c7c3314ef80, C4<1>, C4<1>;
v0x5c7c3300ce70_0 .net "in_a", 0 0, L_0x5c7c3314ef80;  alias, 1 drivers
v0x5c7c3300cf60_0 .net "in_b", 0 0, L_0x5c7c3314ef80;  alias, 1 drivers
v0x5c7c3300d050_0 .net "out", 0 0, L_0x5c7c3314f030;  alias, 1 drivers
S_0x5c7c3300d710 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330097c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3300de40_0 .net "in_a", 0 0, L_0x5c7c3314e9f0;  alias, 1 drivers
v0x5c7c3300dee0_0 .net "out", 0 0, L_0x5c7c3314eaa0;  alias, 1 drivers
S_0x5c7c3300d8e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3300d710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314eaa0 .functor NAND 1, L_0x5c7c3314e9f0, L_0x5c7c3314e9f0, C4<1>, C4<1>;
v0x5c7c3300db50_0 .net "in_a", 0 0, L_0x5c7c3314e9f0;  alias, 1 drivers
v0x5c7c3300dc10_0 .net "in_b", 0 0, L_0x5c7c3314e9f0;  alias, 1 drivers
v0x5c7c3300dd60_0 .net "out", 0 0, L_0x5c7c3314eaa0;  alias, 1 drivers
S_0x5c7c3300dfe0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330097c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3300e7b0_0 .net "in_a", 0 0, L_0x5c7c3314ed10;  alias, 1 drivers
v0x5c7c3300e850_0 .net "out", 0 0, L_0x5c7c3314edc0;  alias, 1 drivers
S_0x5c7c3300e250 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3300dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314edc0 .functor NAND 1, L_0x5c7c3314ed10, L_0x5c7c3314ed10, C4<1>, C4<1>;
v0x5c7c3300e4c0_0 .net "in_a", 0 0, L_0x5c7c3314ed10;  alias, 1 drivers
v0x5c7c3300e580_0 .net "in_b", 0 0, L_0x5c7c3314ed10;  alias, 1 drivers
v0x5c7c3300e6d0_0 .net "out", 0 0, L_0x5c7c3314edc0;  alias, 1 drivers
S_0x5c7c3300e950 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330097c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3300f0f0_0 .net "in_a", 0 0, L_0x5c7c3314f030;  alias, 1 drivers
v0x5c7c3300f190_0 .net "out", 0 0, L_0x5c7c3314f0e0;  alias, 1 drivers
S_0x5c7c3300eb70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3300e950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f0e0 .functor NAND 1, L_0x5c7c3314f030, L_0x5c7c3314f030, C4<1>, C4<1>;
v0x5c7c3300ede0_0 .net "in_a", 0 0, L_0x5c7c3314f030;  alias, 1 drivers
v0x5c7c3300eea0_0 .net "in_b", 0 0, L_0x5c7c3314f030;  alias, 1 drivers
v0x5c7c3300eff0_0 .net "out", 0 0, L_0x5c7c3314f0e0;  alias, 1 drivers
S_0x5c7c33010130 .scope module, "mux_gate3" "Mux" 15 10, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33019490_0 .net "in_a", 0 0, L_0x5c7c331500f0;  1 drivers
v0x5c7c33019530_0 .net "in_b", 0 0, L_0x5c7c33150190;  1 drivers
v0x5c7c33019640_0 .net "out", 0 0, L_0x5c7c3314ff30;  1 drivers
v0x5c7c330196e0_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33019780_0 .net "sel_out", 0 0, L_0x5c7c3314f420;  1 drivers
v0x5c7c33019900_0 .net "temp_a_out", 0 0, L_0x5c7c3314f580;  1 drivers
v0x5c7c33019ab0_0 .net "temp_b_out", 0 0, L_0x5c7c3314f6e0;  1 drivers
S_0x5c7c33010330 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33010130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33011390_0 .net "in_a", 0 0, L_0x5c7c331500f0;  alias, 1 drivers
v0x5c7c33011460_0 .net "in_b", 0 0, L_0x5c7c3314f420;  alias, 1 drivers
v0x5c7c33011530_0 .net "out", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
v0x5c7c33011650_0 .net "temp_out", 0 0, L_0x5c7c3314f4d0;  1 drivers
S_0x5c7c330105a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33010330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f4d0 .functor NAND 1, L_0x5c7c331500f0, L_0x5c7c3314f420, C4<1>, C4<1>;
v0x5c7c33010810_0 .net "in_a", 0 0, L_0x5c7c331500f0;  alias, 1 drivers
v0x5c7c330108f0_0 .net "in_b", 0 0, L_0x5c7c3314f420;  alias, 1 drivers
v0x5c7c330109b0_0 .net "out", 0 0, L_0x5c7c3314f4d0;  alias, 1 drivers
S_0x5c7c33010ad0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33010330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33011210_0 .net "in_a", 0 0, L_0x5c7c3314f4d0;  alias, 1 drivers
v0x5c7c330112b0_0 .net "out", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
S_0x5c7c33010cf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33010ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f580 .functor NAND 1, L_0x5c7c3314f4d0, L_0x5c7c3314f4d0, C4<1>, C4<1>;
v0x5c7c33010f60_0 .net "in_a", 0 0, L_0x5c7c3314f4d0;  alias, 1 drivers
v0x5c7c33011020_0 .net "in_b", 0 0, L_0x5c7c3314f4d0;  alias, 1 drivers
v0x5c7c33011110_0 .net "out", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
S_0x5c7c33011710 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33010130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33012720_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330127c0_0 .net "in_b", 0 0, L_0x5c7c33150190;  alias, 1 drivers
v0x5c7c330128b0_0 .net "out", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
v0x5c7c330129d0_0 .net "temp_out", 0 0, L_0x5c7c3314f630;  1 drivers
S_0x5c7c330118f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33011710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f630 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33150190, C4<1>, C4<1>;
v0x5c7c33011b60_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33011c20_0 .net "in_b", 0 0, L_0x5c7c33150190;  alias, 1 drivers
v0x5c7c33011ce0_0 .net "out", 0 0, L_0x5c7c3314f630;  alias, 1 drivers
S_0x5c7c33011e00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33011710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33012570_0 .net "in_a", 0 0, L_0x5c7c3314f630;  alias, 1 drivers
v0x5c7c33012610_0 .net "out", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
S_0x5c7c33012020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33011e00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f6e0 .functor NAND 1, L_0x5c7c3314f630, L_0x5c7c3314f630, C4<1>, C4<1>;
v0x5c7c33012290_0 .net "in_a", 0 0, L_0x5c7c3314f630;  alias, 1 drivers
v0x5c7c33012380_0 .net "in_b", 0 0, L_0x5c7c3314f630;  alias, 1 drivers
v0x5c7c33012470_0 .net "out", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
S_0x5c7c33012a90 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33010130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33013190_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33013230_0 .net "out", 0 0, L_0x5c7c3314f420;  alias, 1 drivers
S_0x5c7c33012c60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33012a90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f420 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c33012eb0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33012f70_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33013030_0 .net "out", 0 0, L_0x5c7c3314f420;  alias, 1 drivers
S_0x5c7c33013330 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33010130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33018de0_0 .net "branch1_out", 0 0, L_0x5c7c3314f8f0;  1 drivers
v0x5c7c33018f10_0 .net "branch2_out", 0 0, L_0x5c7c3314fc10;  1 drivers
v0x5c7c33019060_0 .net "in_a", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
v0x5c7c33019130_0 .net "in_b", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
v0x5c7c330191d0_0 .net "out", 0 0, L_0x5c7c3314ff30;  alias, 1 drivers
v0x5c7c33019270_0 .net "temp1_out", 0 0, L_0x5c7c3314f840;  1 drivers
v0x5c7c33019310_0 .net "temp2_out", 0 0, L_0x5c7c3314fb60;  1 drivers
v0x5c7c330193b0_0 .net "temp3_out", 0 0, L_0x5c7c3314fe80;  1 drivers
S_0x5c7c33013560 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33013330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33014620_0 .net "in_a", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
v0x5c7c330146c0_0 .net "in_b", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
v0x5c7c33014780_0 .net "out", 0 0, L_0x5c7c3314f840;  alias, 1 drivers
v0x5c7c330148a0_0 .net "temp_out", 0 0, L_0x5c7c3314f790;  1 drivers
S_0x5c7c330137d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33013560;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f790 .functor NAND 1, L_0x5c7c3314f580, L_0x5c7c3314f580, C4<1>, C4<1>;
v0x5c7c33013a40_0 .net "in_a", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
v0x5c7c33013b00_0 .net "in_b", 0 0, L_0x5c7c3314f580;  alias, 1 drivers
v0x5c7c33013c50_0 .net "out", 0 0, L_0x5c7c3314f790;  alias, 1 drivers
S_0x5c7c33013d50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33013560;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33014470_0 .net "in_a", 0 0, L_0x5c7c3314f790;  alias, 1 drivers
v0x5c7c33014510_0 .net "out", 0 0, L_0x5c7c3314f840;  alias, 1 drivers
S_0x5c7c33013f20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33013d50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f840 .functor NAND 1, L_0x5c7c3314f790, L_0x5c7c3314f790, C4<1>, C4<1>;
v0x5c7c33014190_0 .net "in_a", 0 0, L_0x5c7c3314f790;  alias, 1 drivers
v0x5c7c33014280_0 .net "in_b", 0 0, L_0x5c7c3314f790;  alias, 1 drivers
v0x5c7c33014370_0 .net "out", 0 0, L_0x5c7c3314f840;  alias, 1 drivers
S_0x5c7c33014a10 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33013330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33015a40_0 .net "in_a", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
v0x5c7c33015ae0_0 .net "in_b", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
v0x5c7c33015ba0_0 .net "out", 0 0, L_0x5c7c3314fb60;  alias, 1 drivers
v0x5c7c33015cc0_0 .net "temp_out", 0 0, L_0x5c7c3314fab0;  1 drivers
S_0x5c7c33014bf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33014a10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314fab0 .functor NAND 1, L_0x5c7c3314f6e0, L_0x5c7c3314f6e0, C4<1>, C4<1>;
v0x5c7c33014e60_0 .net "in_a", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
v0x5c7c33014f20_0 .net "in_b", 0 0, L_0x5c7c3314f6e0;  alias, 1 drivers
v0x5c7c33015070_0 .net "out", 0 0, L_0x5c7c3314fab0;  alias, 1 drivers
S_0x5c7c33015170 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33014a10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33015890_0 .net "in_a", 0 0, L_0x5c7c3314fab0;  alias, 1 drivers
v0x5c7c33015930_0 .net "out", 0 0, L_0x5c7c3314fb60;  alias, 1 drivers
S_0x5c7c33015340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33015170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314fb60 .functor NAND 1, L_0x5c7c3314fab0, L_0x5c7c3314fab0, C4<1>, C4<1>;
v0x5c7c330155b0_0 .net "in_a", 0 0, L_0x5c7c3314fab0;  alias, 1 drivers
v0x5c7c330156a0_0 .net "in_b", 0 0, L_0x5c7c3314fab0;  alias, 1 drivers
v0x5c7c33015790_0 .net "out", 0 0, L_0x5c7c3314fb60;  alias, 1 drivers
S_0x5c7c33015e30 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33013330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33016e70_0 .net "in_a", 0 0, L_0x5c7c3314f8f0;  alias, 1 drivers
v0x5c7c33016f40_0 .net "in_b", 0 0, L_0x5c7c3314fc10;  alias, 1 drivers
v0x5c7c33017010_0 .net "out", 0 0, L_0x5c7c3314fe80;  alias, 1 drivers
v0x5c7c33017130_0 .net "temp_out", 0 0, L_0x5c7c3314fdd0;  1 drivers
S_0x5c7c33016010 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33015e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314fdd0 .functor NAND 1, L_0x5c7c3314f8f0, L_0x5c7c3314fc10, C4<1>, C4<1>;
v0x5c7c33016260_0 .net "in_a", 0 0, L_0x5c7c3314f8f0;  alias, 1 drivers
v0x5c7c33016340_0 .net "in_b", 0 0, L_0x5c7c3314fc10;  alias, 1 drivers
v0x5c7c33016400_0 .net "out", 0 0, L_0x5c7c3314fdd0;  alias, 1 drivers
S_0x5c7c33016550 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33015e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33016cc0_0 .net "in_a", 0 0, L_0x5c7c3314fdd0;  alias, 1 drivers
v0x5c7c33016d60_0 .net "out", 0 0, L_0x5c7c3314fe80;  alias, 1 drivers
S_0x5c7c33016770 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33016550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314fe80 .functor NAND 1, L_0x5c7c3314fdd0, L_0x5c7c3314fdd0, C4<1>, C4<1>;
v0x5c7c330169e0_0 .net "in_a", 0 0, L_0x5c7c3314fdd0;  alias, 1 drivers
v0x5c7c33016ad0_0 .net "in_b", 0 0, L_0x5c7c3314fdd0;  alias, 1 drivers
v0x5c7c33016bc0_0 .net "out", 0 0, L_0x5c7c3314fe80;  alias, 1 drivers
S_0x5c7c33017280 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33013330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330179b0_0 .net "in_a", 0 0, L_0x5c7c3314f840;  alias, 1 drivers
v0x5c7c33017a50_0 .net "out", 0 0, L_0x5c7c3314f8f0;  alias, 1 drivers
S_0x5c7c33017450 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33017280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314f8f0 .functor NAND 1, L_0x5c7c3314f840, L_0x5c7c3314f840, C4<1>, C4<1>;
v0x5c7c330176c0_0 .net "in_a", 0 0, L_0x5c7c3314f840;  alias, 1 drivers
v0x5c7c33017780_0 .net "in_b", 0 0, L_0x5c7c3314f840;  alias, 1 drivers
v0x5c7c330178d0_0 .net "out", 0 0, L_0x5c7c3314f8f0;  alias, 1 drivers
S_0x5c7c33017b50 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33013330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33018320_0 .net "in_a", 0 0, L_0x5c7c3314fb60;  alias, 1 drivers
v0x5c7c330183c0_0 .net "out", 0 0, L_0x5c7c3314fc10;  alias, 1 drivers
S_0x5c7c33017dc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33017b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314fc10 .functor NAND 1, L_0x5c7c3314fb60, L_0x5c7c3314fb60, C4<1>, C4<1>;
v0x5c7c33018030_0 .net "in_a", 0 0, L_0x5c7c3314fb60;  alias, 1 drivers
v0x5c7c330180f0_0 .net "in_b", 0 0, L_0x5c7c3314fb60;  alias, 1 drivers
v0x5c7c33018240_0 .net "out", 0 0, L_0x5c7c3314fc10;  alias, 1 drivers
S_0x5c7c330184c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33013330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33018c60_0 .net "in_a", 0 0, L_0x5c7c3314fe80;  alias, 1 drivers
v0x5c7c33018d00_0 .net "out", 0 0, L_0x5c7c3314ff30;  alias, 1 drivers
S_0x5c7c330186e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330184c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3314ff30 .functor NAND 1, L_0x5c7c3314fe80, L_0x5c7c3314fe80, C4<1>, C4<1>;
v0x5c7c33018950_0 .net "in_a", 0 0, L_0x5c7c3314fe80;  alias, 1 drivers
v0x5c7c33018a10_0 .net "in_b", 0 0, L_0x5c7c3314fe80;  alias, 1 drivers
v0x5c7c33018b60_0 .net "out", 0 0, L_0x5c7c3314ff30;  alias, 1 drivers
S_0x5c7c33019ca0 .scope module, "mux_gate4" "Mux" 15 11, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33023810_0 .net "in_a", 0 0, L_0x5c7c33150f00;  1 drivers
v0x5c7c330238b0_0 .net "in_b", 0 0, L_0x5c7c33150fa0;  1 drivers
v0x5c7c330239c0_0 .net "out", 0 0, L_0x5c7c33150d40;  1 drivers
v0x5c7c33023a60_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33023b00_0 .net "sel_out", 0 0, L_0x5c7c33150230;  1 drivers
v0x5c7c33023c80_0 .net "temp_a_out", 0 0, L_0x5c7c33150390;  1 drivers
v0x5c7c33023e30_0 .net "temp_b_out", 0 0, L_0x5c7c331504f0;  1 drivers
S_0x5c7c33019ea0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33019ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3301af00_0 .net "in_a", 0 0, L_0x5c7c33150f00;  alias, 1 drivers
v0x5c7c3301afd0_0 .net "in_b", 0 0, L_0x5c7c33150230;  alias, 1 drivers
v0x5c7c3301b0a0_0 .net "out", 0 0, L_0x5c7c33150390;  alias, 1 drivers
v0x5c7c3301b1c0_0 .net "temp_out", 0 0, L_0x5c7c331502e0;  1 drivers
S_0x5c7c3301a110 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33019ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331502e0 .functor NAND 1, L_0x5c7c33150f00, L_0x5c7c33150230, C4<1>, C4<1>;
v0x5c7c3301a380_0 .net "in_a", 0 0, L_0x5c7c33150f00;  alias, 1 drivers
v0x5c7c3301a460_0 .net "in_b", 0 0, L_0x5c7c33150230;  alias, 1 drivers
v0x5c7c3301a520_0 .net "out", 0 0, L_0x5c7c331502e0;  alias, 1 drivers
S_0x5c7c3301a640 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33019ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3301ad80_0 .net "in_a", 0 0, L_0x5c7c331502e0;  alias, 1 drivers
v0x5c7c3301ae20_0 .net "out", 0 0, L_0x5c7c33150390;  alias, 1 drivers
S_0x5c7c3301a860 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3301a640;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150390 .functor NAND 1, L_0x5c7c331502e0, L_0x5c7c331502e0, C4<1>, C4<1>;
v0x5c7c3301aad0_0 .net "in_a", 0 0, L_0x5c7c331502e0;  alias, 1 drivers
v0x5c7c3301ab90_0 .net "in_b", 0 0, L_0x5c7c331502e0;  alias, 1 drivers
v0x5c7c3301ac80_0 .net "out", 0 0, L_0x5c7c33150390;  alias, 1 drivers
S_0x5c7c3301b280 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33019ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3301c290_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3301c330_0 .net "in_b", 0 0, L_0x5c7c33150fa0;  alias, 1 drivers
v0x5c7c3301c420_0 .net "out", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
v0x5c7c3301c540_0 .net "temp_out", 0 0, L_0x5c7c33150440;  1 drivers
S_0x5c7c3301b460 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3301b280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150440 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33150fa0, C4<1>, C4<1>;
v0x5c7c3301b6d0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3301b790_0 .net "in_b", 0 0, L_0x5c7c33150fa0;  alias, 1 drivers
v0x5c7c3301b850_0 .net "out", 0 0, L_0x5c7c33150440;  alias, 1 drivers
S_0x5c7c3301b970 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3301b280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3301c0e0_0 .net "in_a", 0 0, L_0x5c7c33150440;  alias, 1 drivers
v0x5c7c3301c180_0 .net "out", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
S_0x5c7c3301bb90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3301b970;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331504f0 .functor NAND 1, L_0x5c7c33150440, L_0x5c7c33150440, C4<1>, C4<1>;
v0x5c7c3301be00_0 .net "in_a", 0 0, L_0x5c7c33150440;  alias, 1 drivers
v0x5c7c3301bef0_0 .net "in_b", 0 0, L_0x5c7c33150440;  alias, 1 drivers
v0x5c7c3301bfe0_0 .net "out", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
S_0x5c7c3301c600 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33019ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3301cd00_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3301d5b0_0 .net "out", 0 0, L_0x5c7c33150230;  alias, 1 drivers
S_0x5c7c3301c7d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3301c600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150230 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c3301ca20_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3301cae0_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3301cba0_0 .net "out", 0 0, L_0x5c7c33150230;  alias, 1 drivers
S_0x5c7c3301d6b0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33019ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33023160_0 .net "branch1_out", 0 0, L_0x5c7c33150700;  1 drivers
v0x5c7c33023290_0 .net "branch2_out", 0 0, L_0x5c7c33150a20;  1 drivers
v0x5c7c330233e0_0 .net "in_a", 0 0, L_0x5c7c33150390;  alias, 1 drivers
v0x5c7c330234b0_0 .net "in_b", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
v0x5c7c33023550_0 .net "out", 0 0, L_0x5c7c33150d40;  alias, 1 drivers
v0x5c7c330235f0_0 .net "temp1_out", 0 0, L_0x5c7c33150650;  1 drivers
v0x5c7c33023690_0 .net "temp2_out", 0 0, L_0x5c7c33150970;  1 drivers
v0x5c7c33023730_0 .net "temp3_out", 0 0, L_0x5c7c33150c90;  1 drivers
S_0x5c7c3301d8e0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c3301d6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3301e9a0_0 .net "in_a", 0 0, L_0x5c7c33150390;  alias, 1 drivers
v0x5c7c3301ea40_0 .net "in_b", 0 0, L_0x5c7c33150390;  alias, 1 drivers
v0x5c7c3301eb00_0 .net "out", 0 0, L_0x5c7c33150650;  alias, 1 drivers
v0x5c7c3301ec20_0 .net "temp_out", 0 0, L_0x5c7c331505a0;  1 drivers
S_0x5c7c3301db50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3301d8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331505a0 .functor NAND 1, L_0x5c7c33150390, L_0x5c7c33150390, C4<1>, C4<1>;
v0x5c7c3301ddc0_0 .net "in_a", 0 0, L_0x5c7c33150390;  alias, 1 drivers
v0x5c7c3301de80_0 .net "in_b", 0 0, L_0x5c7c33150390;  alias, 1 drivers
v0x5c7c3301dfd0_0 .net "out", 0 0, L_0x5c7c331505a0;  alias, 1 drivers
S_0x5c7c3301e0d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3301d8e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3301e7f0_0 .net "in_a", 0 0, L_0x5c7c331505a0;  alias, 1 drivers
v0x5c7c3301e890_0 .net "out", 0 0, L_0x5c7c33150650;  alias, 1 drivers
S_0x5c7c3301e2a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3301e0d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150650 .functor NAND 1, L_0x5c7c331505a0, L_0x5c7c331505a0, C4<1>, C4<1>;
v0x5c7c3301e510_0 .net "in_a", 0 0, L_0x5c7c331505a0;  alias, 1 drivers
v0x5c7c3301e600_0 .net "in_b", 0 0, L_0x5c7c331505a0;  alias, 1 drivers
v0x5c7c3301e6f0_0 .net "out", 0 0, L_0x5c7c33150650;  alias, 1 drivers
S_0x5c7c3301ed90 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c3301d6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3301fdc0_0 .net "in_a", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
v0x5c7c3301fe60_0 .net "in_b", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
v0x5c7c3301ff20_0 .net "out", 0 0, L_0x5c7c33150970;  alias, 1 drivers
v0x5c7c33020040_0 .net "temp_out", 0 0, L_0x5c7c331508c0;  1 drivers
S_0x5c7c3301ef70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3301ed90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331508c0 .functor NAND 1, L_0x5c7c331504f0, L_0x5c7c331504f0, C4<1>, C4<1>;
v0x5c7c3301f1e0_0 .net "in_a", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
v0x5c7c3301f2a0_0 .net "in_b", 0 0, L_0x5c7c331504f0;  alias, 1 drivers
v0x5c7c3301f3f0_0 .net "out", 0 0, L_0x5c7c331508c0;  alias, 1 drivers
S_0x5c7c3301f4f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3301ed90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3301fc10_0 .net "in_a", 0 0, L_0x5c7c331508c0;  alias, 1 drivers
v0x5c7c3301fcb0_0 .net "out", 0 0, L_0x5c7c33150970;  alias, 1 drivers
S_0x5c7c3301f6c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3301f4f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150970 .functor NAND 1, L_0x5c7c331508c0, L_0x5c7c331508c0, C4<1>, C4<1>;
v0x5c7c3301f930_0 .net "in_a", 0 0, L_0x5c7c331508c0;  alias, 1 drivers
v0x5c7c3301fa20_0 .net "in_b", 0 0, L_0x5c7c331508c0;  alias, 1 drivers
v0x5c7c3301fb10_0 .net "out", 0 0, L_0x5c7c33150970;  alias, 1 drivers
S_0x5c7c330201b0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c3301d6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330211f0_0 .net "in_a", 0 0, L_0x5c7c33150700;  alias, 1 drivers
v0x5c7c330212c0_0 .net "in_b", 0 0, L_0x5c7c33150a20;  alias, 1 drivers
v0x5c7c33021390_0 .net "out", 0 0, L_0x5c7c33150c90;  alias, 1 drivers
v0x5c7c330214b0_0 .net "temp_out", 0 0, L_0x5c7c33150be0;  1 drivers
S_0x5c7c33020390 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330201b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150be0 .functor NAND 1, L_0x5c7c33150700, L_0x5c7c33150a20, C4<1>, C4<1>;
v0x5c7c330205e0_0 .net "in_a", 0 0, L_0x5c7c33150700;  alias, 1 drivers
v0x5c7c330206c0_0 .net "in_b", 0 0, L_0x5c7c33150a20;  alias, 1 drivers
v0x5c7c33020780_0 .net "out", 0 0, L_0x5c7c33150be0;  alias, 1 drivers
S_0x5c7c330208d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330201b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33021040_0 .net "in_a", 0 0, L_0x5c7c33150be0;  alias, 1 drivers
v0x5c7c330210e0_0 .net "out", 0 0, L_0x5c7c33150c90;  alias, 1 drivers
S_0x5c7c33020af0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330208d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150c90 .functor NAND 1, L_0x5c7c33150be0, L_0x5c7c33150be0, C4<1>, C4<1>;
v0x5c7c33020d60_0 .net "in_a", 0 0, L_0x5c7c33150be0;  alias, 1 drivers
v0x5c7c33020e50_0 .net "in_b", 0 0, L_0x5c7c33150be0;  alias, 1 drivers
v0x5c7c33020f40_0 .net "out", 0 0, L_0x5c7c33150c90;  alias, 1 drivers
S_0x5c7c33021600 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c3301d6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33021d30_0 .net "in_a", 0 0, L_0x5c7c33150650;  alias, 1 drivers
v0x5c7c33021dd0_0 .net "out", 0 0, L_0x5c7c33150700;  alias, 1 drivers
S_0x5c7c330217d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33021600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150700 .functor NAND 1, L_0x5c7c33150650, L_0x5c7c33150650, C4<1>, C4<1>;
v0x5c7c33021a40_0 .net "in_a", 0 0, L_0x5c7c33150650;  alias, 1 drivers
v0x5c7c33021b00_0 .net "in_b", 0 0, L_0x5c7c33150650;  alias, 1 drivers
v0x5c7c33021c50_0 .net "out", 0 0, L_0x5c7c33150700;  alias, 1 drivers
S_0x5c7c33021ed0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c3301d6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330226a0_0 .net "in_a", 0 0, L_0x5c7c33150970;  alias, 1 drivers
v0x5c7c33022740_0 .net "out", 0 0, L_0x5c7c33150a20;  alias, 1 drivers
S_0x5c7c33022140 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33021ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150a20 .functor NAND 1, L_0x5c7c33150970, L_0x5c7c33150970, C4<1>, C4<1>;
v0x5c7c330223b0_0 .net "in_a", 0 0, L_0x5c7c33150970;  alias, 1 drivers
v0x5c7c33022470_0 .net "in_b", 0 0, L_0x5c7c33150970;  alias, 1 drivers
v0x5c7c330225c0_0 .net "out", 0 0, L_0x5c7c33150a20;  alias, 1 drivers
S_0x5c7c33022840 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c3301d6b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33022fe0_0 .net "in_a", 0 0, L_0x5c7c33150c90;  alias, 1 drivers
v0x5c7c33023080_0 .net "out", 0 0, L_0x5c7c33150d40;  alias, 1 drivers
S_0x5c7c33022a60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33022840;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33150d40 .functor NAND 1, L_0x5c7c33150c90, L_0x5c7c33150c90, C4<1>, C4<1>;
v0x5c7c33022cd0_0 .net "in_a", 0 0, L_0x5c7c33150c90;  alias, 1 drivers
v0x5c7c33022d90_0 .net "in_b", 0 0, L_0x5c7c33150c90;  alias, 1 drivers
v0x5c7c33022ee0_0 .net "out", 0 0, L_0x5c7c33150d40;  alias, 1 drivers
S_0x5c7c33024020 .scope module, "mux_gate5" "Mux" 15 12, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c3302d380_0 .net "in_a", 0 0, L_0x5c7c33151d70;  1 drivers
v0x5c7c3302d420_0 .net "in_b", 0 0, L_0x5c7c33151e10;  1 drivers
v0x5c7c3302d530_0 .net "out", 0 0, L_0x5c7c33151bb0;  1 drivers
v0x5c7c3302d5d0_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3302d670_0 .net "sel_out", 0 0, L_0x5c7c331510a0;  1 drivers
v0x5c7c3302d7f0_0 .net "temp_a_out", 0 0, L_0x5c7c33151200;  1 drivers
v0x5c7c3302d9a0_0 .net "temp_b_out", 0 0, L_0x5c7c33151360;  1 drivers
S_0x5c7c33024220 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33024020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33025280_0 .net "in_a", 0 0, L_0x5c7c33151d70;  alias, 1 drivers
v0x5c7c33025350_0 .net "in_b", 0 0, L_0x5c7c331510a0;  alias, 1 drivers
v0x5c7c33025420_0 .net "out", 0 0, L_0x5c7c33151200;  alias, 1 drivers
v0x5c7c33025540_0 .net "temp_out", 0 0, L_0x5c7c33151150;  1 drivers
S_0x5c7c33024490 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33024220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151150 .functor NAND 1, L_0x5c7c33151d70, L_0x5c7c331510a0, C4<1>, C4<1>;
v0x5c7c33024700_0 .net "in_a", 0 0, L_0x5c7c33151d70;  alias, 1 drivers
v0x5c7c330247e0_0 .net "in_b", 0 0, L_0x5c7c331510a0;  alias, 1 drivers
v0x5c7c330248a0_0 .net "out", 0 0, L_0x5c7c33151150;  alias, 1 drivers
S_0x5c7c330249c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33024220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33025100_0 .net "in_a", 0 0, L_0x5c7c33151150;  alias, 1 drivers
v0x5c7c330251a0_0 .net "out", 0 0, L_0x5c7c33151200;  alias, 1 drivers
S_0x5c7c33024be0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330249c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151200 .functor NAND 1, L_0x5c7c33151150, L_0x5c7c33151150, C4<1>, C4<1>;
v0x5c7c33024e50_0 .net "in_a", 0 0, L_0x5c7c33151150;  alias, 1 drivers
v0x5c7c33024f10_0 .net "in_b", 0 0, L_0x5c7c33151150;  alias, 1 drivers
v0x5c7c33025000_0 .net "out", 0 0, L_0x5c7c33151200;  alias, 1 drivers
S_0x5c7c33025600 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33024020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33026610_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330266b0_0 .net "in_b", 0 0, L_0x5c7c33151e10;  alias, 1 drivers
v0x5c7c330267a0_0 .net "out", 0 0, L_0x5c7c33151360;  alias, 1 drivers
v0x5c7c330268c0_0 .net "temp_out", 0 0, L_0x5c7c331512b0;  1 drivers
S_0x5c7c330257e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33025600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331512b0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33151e10, C4<1>, C4<1>;
v0x5c7c33025a50_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33025b10_0 .net "in_b", 0 0, L_0x5c7c33151e10;  alias, 1 drivers
v0x5c7c33025bd0_0 .net "out", 0 0, L_0x5c7c331512b0;  alias, 1 drivers
S_0x5c7c33025cf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33025600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33026460_0 .net "in_a", 0 0, L_0x5c7c331512b0;  alias, 1 drivers
v0x5c7c33026500_0 .net "out", 0 0, L_0x5c7c33151360;  alias, 1 drivers
S_0x5c7c33025f10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33025cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151360 .functor NAND 1, L_0x5c7c331512b0, L_0x5c7c331512b0, C4<1>, C4<1>;
v0x5c7c33026180_0 .net "in_a", 0 0, L_0x5c7c331512b0;  alias, 1 drivers
v0x5c7c33026270_0 .net "in_b", 0 0, L_0x5c7c331512b0;  alias, 1 drivers
v0x5c7c33026360_0 .net "out", 0 0, L_0x5c7c33151360;  alias, 1 drivers
S_0x5c7c33026980 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33024020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33027080_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33027120_0 .net "out", 0 0, L_0x5c7c331510a0;  alias, 1 drivers
S_0x5c7c33026b50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33026980;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331510a0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c33026da0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33026e60_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33026f20_0 .net "out", 0 0, L_0x5c7c331510a0;  alias, 1 drivers
S_0x5c7c33027220 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33024020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3302ccd0_0 .net "branch1_out", 0 0, L_0x5c7c33151570;  1 drivers
v0x5c7c3302ce00_0 .net "branch2_out", 0 0, L_0x5c7c33151890;  1 drivers
v0x5c7c3302cf50_0 .net "in_a", 0 0, L_0x5c7c33151200;  alias, 1 drivers
v0x5c7c3302d020_0 .net "in_b", 0 0, L_0x5c7c33151360;  alias, 1 drivers
v0x5c7c3302d0c0_0 .net "out", 0 0, L_0x5c7c33151bb0;  alias, 1 drivers
v0x5c7c3302d160_0 .net "temp1_out", 0 0, L_0x5c7c331514c0;  1 drivers
v0x5c7c3302d200_0 .net "temp2_out", 0 0, L_0x5c7c331517e0;  1 drivers
v0x5c7c3302d2a0_0 .net "temp3_out", 0 0, L_0x5c7c33151b00;  1 drivers
S_0x5c7c33027450 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33027220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33028510_0 .net "in_a", 0 0, L_0x5c7c33151200;  alias, 1 drivers
v0x5c7c330285b0_0 .net "in_b", 0 0, L_0x5c7c33151200;  alias, 1 drivers
v0x5c7c33028670_0 .net "out", 0 0, L_0x5c7c331514c0;  alias, 1 drivers
v0x5c7c33028790_0 .net "temp_out", 0 0, L_0x5c7c33151410;  1 drivers
S_0x5c7c330276c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33027450;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151410 .functor NAND 1, L_0x5c7c33151200, L_0x5c7c33151200, C4<1>, C4<1>;
v0x5c7c33027930_0 .net "in_a", 0 0, L_0x5c7c33151200;  alias, 1 drivers
v0x5c7c330279f0_0 .net "in_b", 0 0, L_0x5c7c33151200;  alias, 1 drivers
v0x5c7c33027b40_0 .net "out", 0 0, L_0x5c7c33151410;  alias, 1 drivers
S_0x5c7c33027c40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33027450;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33028360_0 .net "in_a", 0 0, L_0x5c7c33151410;  alias, 1 drivers
v0x5c7c33028400_0 .net "out", 0 0, L_0x5c7c331514c0;  alias, 1 drivers
S_0x5c7c33027e10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33027c40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331514c0 .functor NAND 1, L_0x5c7c33151410, L_0x5c7c33151410, C4<1>, C4<1>;
v0x5c7c33028080_0 .net "in_a", 0 0, L_0x5c7c33151410;  alias, 1 drivers
v0x5c7c33028170_0 .net "in_b", 0 0, L_0x5c7c33151410;  alias, 1 drivers
v0x5c7c33028260_0 .net "out", 0 0, L_0x5c7c331514c0;  alias, 1 drivers
S_0x5c7c33028900 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33027220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33029930_0 .net "in_a", 0 0, L_0x5c7c33151360;  alias, 1 drivers
v0x5c7c330299d0_0 .net "in_b", 0 0, L_0x5c7c33151360;  alias, 1 drivers
v0x5c7c33029a90_0 .net "out", 0 0, L_0x5c7c331517e0;  alias, 1 drivers
v0x5c7c33029bb0_0 .net "temp_out", 0 0, L_0x5c7c33151730;  1 drivers
S_0x5c7c33028ae0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33028900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151730 .functor NAND 1, L_0x5c7c33151360, L_0x5c7c33151360, C4<1>, C4<1>;
v0x5c7c33028d50_0 .net "in_a", 0 0, L_0x5c7c33151360;  alias, 1 drivers
v0x5c7c33028e10_0 .net "in_b", 0 0, L_0x5c7c33151360;  alias, 1 drivers
v0x5c7c33028f60_0 .net "out", 0 0, L_0x5c7c33151730;  alias, 1 drivers
S_0x5c7c33029060 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33028900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33029780_0 .net "in_a", 0 0, L_0x5c7c33151730;  alias, 1 drivers
v0x5c7c33029820_0 .net "out", 0 0, L_0x5c7c331517e0;  alias, 1 drivers
S_0x5c7c33029230 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33029060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331517e0 .functor NAND 1, L_0x5c7c33151730, L_0x5c7c33151730, C4<1>, C4<1>;
v0x5c7c330294a0_0 .net "in_a", 0 0, L_0x5c7c33151730;  alias, 1 drivers
v0x5c7c33029590_0 .net "in_b", 0 0, L_0x5c7c33151730;  alias, 1 drivers
v0x5c7c33029680_0 .net "out", 0 0, L_0x5c7c331517e0;  alias, 1 drivers
S_0x5c7c33029d20 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33027220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3302ad60_0 .net "in_a", 0 0, L_0x5c7c33151570;  alias, 1 drivers
v0x5c7c3302ae30_0 .net "in_b", 0 0, L_0x5c7c33151890;  alias, 1 drivers
v0x5c7c3302af00_0 .net "out", 0 0, L_0x5c7c33151b00;  alias, 1 drivers
v0x5c7c3302b020_0 .net "temp_out", 0 0, L_0x5c7c33151a50;  1 drivers
S_0x5c7c33029f00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33029d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151a50 .functor NAND 1, L_0x5c7c33151570, L_0x5c7c33151890, C4<1>, C4<1>;
v0x5c7c3302a150_0 .net "in_a", 0 0, L_0x5c7c33151570;  alias, 1 drivers
v0x5c7c3302a230_0 .net "in_b", 0 0, L_0x5c7c33151890;  alias, 1 drivers
v0x5c7c3302a2f0_0 .net "out", 0 0, L_0x5c7c33151a50;  alias, 1 drivers
S_0x5c7c3302a440 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33029d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3302abb0_0 .net "in_a", 0 0, L_0x5c7c33151a50;  alias, 1 drivers
v0x5c7c3302ac50_0 .net "out", 0 0, L_0x5c7c33151b00;  alias, 1 drivers
S_0x5c7c3302a660 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3302a440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151b00 .functor NAND 1, L_0x5c7c33151a50, L_0x5c7c33151a50, C4<1>, C4<1>;
v0x5c7c3302a8d0_0 .net "in_a", 0 0, L_0x5c7c33151a50;  alias, 1 drivers
v0x5c7c3302a9c0_0 .net "in_b", 0 0, L_0x5c7c33151a50;  alias, 1 drivers
v0x5c7c3302aab0_0 .net "out", 0 0, L_0x5c7c33151b00;  alias, 1 drivers
S_0x5c7c3302b170 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33027220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3302b8a0_0 .net "in_a", 0 0, L_0x5c7c331514c0;  alias, 1 drivers
v0x5c7c3302b940_0 .net "out", 0 0, L_0x5c7c33151570;  alias, 1 drivers
S_0x5c7c3302b340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3302b170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151570 .functor NAND 1, L_0x5c7c331514c0, L_0x5c7c331514c0, C4<1>, C4<1>;
v0x5c7c3302b5b0_0 .net "in_a", 0 0, L_0x5c7c331514c0;  alias, 1 drivers
v0x5c7c3302b670_0 .net "in_b", 0 0, L_0x5c7c331514c0;  alias, 1 drivers
v0x5c7c3302b7c0_0 .net "out", 0 0, L_0x5c7c33151570;  alias, 1 drivers
S_0x5c7c3302ba40 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33027220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3302c210_0 .net "in_a", 0 0, L_0x5c7c331517e0;  alias, 1 drivers
v0x5c7c3302c2b0_0 .net "out", 0 0, L_0x5c7c33151890;  alias, 1 drivers
S_0x5c7c3302bcb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3302ba40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151890 .functor NAND 1, L_0x5c7c331517e0, L_0x5c7c331517e0, C4<1>, C4<1>;
v0x5c7c3302bf20_0 .net "in_a", 0 0, L_0x5c7c331517e0;  alias, 1 drivers
v0x5c7c3302bfe0_0 .net "in_b", 0 0, L_0x5c7c331517e0;  alias, 1 drivers
v0x5c7c3302c130_0 .net "out", 0 0, L_0x5c7c33151890;  alias, 1 drivers
S_0x5c7c3302c3b0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33027220;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3302cb50_0 .net "in_a", 0 0, L_0x5c7c33151b00;  alias, 1 drivers
v0x5c7c3302cbf0_0 .net "out", 0 0, L_0x5c7c33151bb0;  alias, 1 drivers
S_0x5c7c3302c5d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3302c3b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151bb0 .functor NAND 1, L_0x5c7c33151b00, L_0x5c7c33151b00, C4<1>, C4<1>;
v0x5c7c3302c840_0 .net "in_a", 0 0, L_0x5c7c33151b00;  alias, 1 drivers
v0x5c7c3302c900_0 .net "in_b", 0 0, L_0x5c7c33151b00;  alias, 1 drivers
v0x5c7c3302ca50_0 .net "out", 0 0, L_0x5c7c33151bb0;  alias, 1 drivers
S_0x5c7c3302db90 .scope module, "mux_gate6" "Mux" 15 13, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33036ef0_0 .net "in_a", 0 0, L_0x5c7c33152bf0;  1 drivers
v0x5c7c33036f90_0 .net "in_b", 0 0, L_0x5c7c33152da0;  1 drivers
v0x5c7c330370a0_0 .net "out", 0 0, L_0x5c7c33152a30;  1 drivers
v0x5c7c33037140_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330371e0_0 .net "sel_out", 0 0, L_0x5c7c33151f20;  1 drivers
v0x5c7c33037360_0 .net "temp_a_out", 0 0, L_0x5c7c33152080;  1 drivers
v0x5c7c33037510_0 .net "temp_b_out", 0 0, L_0x5c7c331521e0;  1 drivers
S_0x5c7c3302dd90 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c3302db90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3302edf0_0 .net "in_a", 0 0, L_0x5c7c33152bf0;  alias, 1 drivers
v0x5c7c3302eec0_0 .net "in_b", 0 0, L_0x5c7c33151f20;  alias, 1 drivers
v0x5c7c3302ef90_0 .net "out", 0 0, L_0x5c7c33152080;  alias, 1 drivers
v0x5c7c3302f0b0_0 .net "temp_out", 0 0, L_0x5c7c33151fd0;  1 drivers
S_0x5c7c3302e000 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3302dd90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151fd0 .functor NAND 1, L_0x5c7c33152bf0, L_0x5c7c33151f20, C4<1>, C4<1>;
v0x5c7c3302e270_0 .net "in_a", 0 0, L_0x5c7c33152bf0;  alias, 1 drivers
v0x5c7c3302e350_0 .net "in_b", 0 0, L_0x5c7c33151f20;  alias, 1 drivers
v0x5c7c3302e410_0 .net "out", 0 0, L_0x5c7c33151fd0;  alias, 1 drivers
S_0x5c7c3302e530 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3302dd90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3302ec70_0 .net "in_a", 0 0, L_0x5c7c33151fd0;  alias, 1 drivers
v0x5c7c3302ed10_0 .net "out", 0 0, L_0x5c7c33152080;  alias, 1 drivers
S_0x5c7c3302e750 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3302e530;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152080 .functor NAND 1, L_0x5c7c33151fd0, L_0x5c7c33151fd0, C4<1>, C4<1>;
v0x5c7c3302e9c0_0 .net "in_a", 0 0, L_0x5c7c33151fd0;  alias, 1 drivers
v0x5c7c3302ea80_0 .net "in_b", 0 0, L_0x5c7c33151fd0;  alias, 1 drivers
v0x5c7c3302eb70_0 .net "out", 0 0, L_0x5c7c33152080;  alias, 1 drivers
S_0x5c7c3302f170 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c3302db90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33030180_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33030220_0 .net "in_b", 0 0, L_0x5c7c33152da0;  alias, 1 drivers
v0x5c7c33030310_0 .net "out", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
v0x5c7c33030430_0 .net "temp_out", 0 0, L_0x5c7c33152130;  1 drivers
S_0x5c7c3302f350 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3302f170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152130 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33152da0, C4<1>, C4<1>;
v0x5c7c3302f5c0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3302f680_0 .net "in_b", 0 0, L_0x5c7c33152da0;  alias, 1 drivers
v0x5c7c3302f740_0 .net "out", 0 0, L_0x5c7c33152130;  alias, 1 drivers
S_0x5c7c3302f860 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3302f170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3302ffd0_0 .net "in_a", 0 0, L_0x5c7c33152130;  alias, 1 drivers
v0x5c7c33030070_0 .net "out", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
S_0x5c7c3302fa80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3302f860;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331521e0 .functor NAND 1, L_0x5c7c33152130, L_0x5c7c33152130, C4<1>, C4<1>;
v0x5c7c3302fcf0_0 .net "in_a", 0 0, L_0x5c7c33152130;  alias, 1 drivers
v0x5c7c3302fde0_0 .net "in_b", 0 0, L_0x5c7c33152130;  alias, 1 drivers
v0x5c7c3302fed0_0 .net "out", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
S_0x5c7c330304f0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c3302db90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33030bf0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33030c90_0 .net "out", 0 0, L_0x5c7c33151f20;  alias, 1 drivers
S_0x5c7c330306c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330304f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151f20 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c33030910_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330309d0_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33030a90_0 .net "out", 0 0, L_0x5c7c33151f20;  alias, 1 drivers
S_0x5c7c33030d90 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c3302db90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33036840_0 .net "branch1_out", 0 0, L_0x5c7c331523f0;  1 drivers
v0x5c7c33036970_0 .net "branch2_out", 0 0, L_0x5c7c33152710;  1 drivers
v0x5c7c33036ac0_0 .net "in_a", 0 0, L_0x5c7c33152080;  alias, 1 drivers
v0x5c7c33036b90_0 .net "in_b", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
v0x5c7c33036c30_0 .net "out", 0 0, L_0x5c7c33152a30;  alias, 1 drivers
v0x5c7c33036cd0_0 .net "temp1_out", 0 0, L_0x5c7c33152340;  1 drivers
v0x5c7c33036d70_0 .net "temp2_out", 0 0, L_0x5c7c33152660;  1 drivers
v0x5c7c33036e10_0 .net "temp3_out", 0 0, L_0x5c7c33152980;  1 drivers
S_0x5c7c33030fc0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33030d90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33032080_0 .net "in_a", 0 0, L_0x5c7c33152080;  alias, 1 drivers
v0x5c7c33032120_0 .net "in_b", 0 0, L_0x5c7c33152080;  alias, 1 drivers
v0x5c7c330321e0_0 .net "out", 0 0, L_0x5c7c33152340;  alias, 1 drivers
v0x5c7c33032300_0 .net "temp_out", 0 0, L_0x5c7c33152290;  1 drivers
S_0x5c7c33031230 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33030fc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152290 .functor NAND 1, L_0x5c7c33152080, L_0x5c7c33152080, C4<1>, C4<1>;
v0x5c7c330314a0_0 .net "in_a", 0 0, L_0x5c7c33152080;  alias, 1 drivers
v0x5c7c33031560_0 .net "in_b", 0 0, L_0x5c7c33152080;  alias, 1 drivers
v0x5c7c330316b0_0 .net "out", 0 0, L_0x5c7c33152290;  alias, 1 drivers
S_0x5c7c330317b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33030fc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33031ed0_0 .net "in_a", 0 0, L_0x5c7c33152290;  alias, 1 drivers
v0x5c7c33031f70_0 .net "out", 0 0, L_0x5c7c33152340;  alias, 1 drivers
S_0x5c7c33031980 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330317b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152340 .functor NAND 1, L_0x5c7c33152290, L_0x5c7c33152290, C4<1>, C4<1>;
v0x5c7c33031bf0_0 .net "in_a", 0 0, L_0x5c7c33152290;  alias, 1 drivers
v0x5c7c33031ce0_0 .net "in_b", 0 0, L_0x5c7c33152290;  alias, 1 drivers
v0x5c7c33031dd0_0 .net "out", 0 0, L_0x5c7c33152340;  alias, 1 drivers
S_0x5c7c33032470 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33030d90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330334a0_0 .net "in_a", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
v0x5c7c33033540_0 .net "in_b", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
v0x5c7c33033600_0 .net "out", 0 0, L_0x5c7c33152660;  alias, 1 drivers
v0x5c7c33033720_0 .net "temp_out", 0 0, L_0x5c7c331525b0;  1 drivers
S_0x5c7c33032650 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33032470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331525b0 .functor NAND 1, L_0x5c7c331521e0, L_0x5c7c331521e0, C4<1>, C4<1>;
v0x5c7c330328c0_0 .net "in_a", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
v0x5c7c33032980_0 .net "in_b", 0 0, L_0x5c7c331521e0;  alias, 1 drivers
v0x5c7c33032ad0_0 .net "out", 0 0, L_0x5c7c331525b0;  alias, 1 drivers
S_0x5c7c33032bd0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33032470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330332f0_0 .net "in_a", 0 0, L_0x5c7c331525b0;  alias, 1 drivers
v0x5c7c33033390_0 .net "out", 0 0, L_0x5c7c33152660;  alias, 1 drivers
S_0x5c7c33032da0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33032bd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152660 .functor NAND 1, L_0x5c7c331525b0, L_0x5c7c331525b0, C4<1>, C4<1>;
v0x5c7c33033010_0 .net "in_a", 0 0, L_0x5c7c331525b0;  alias, 1 drivers
v0x5c7c33033100_0 .net "in_b", 0 0, L_0x5c7c331525b0;  alias, 1 drivers
v0x5c7c330331f0_0 .net "out", 0 0, L_0x5c7c33152660;  alias, 1 drivers
S_0x5c7c33033890 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33030d90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330348d0_0 .net "in_a", 0 0, L_0x5c7c331523f0;  alias, 1 drivers
v0x5c7c330349a0_0 .net "in_b", 0 0, L_0x5c7c33152710;  alias, 1 drivers
v0x5c7c33034a70_0 .net "out", 0 0, L_0x5c7c33152980;  alias, 1 drivers
v0x5c7c33034b90_0 .net "temp_out", 0 0, L_0x5c7c331528d0;  1 drivers
S_0x5c7c33033a70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33033890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331528d0 .functor NAND 1, L_0x5c7c331523f0, L_0x5c7c33152710, C4<1>, C4<1>;
v0x5c7c33033cc0_0 .net "in_a", 0 0, L_0x5c7c331523f0;  alias, 1 drivers
v0x5c7c33033da0_0 .net "in_b", 0 0, L_0x5c7c33152710;  alias, 1 drivers
v0x5c7c33033e60_0 .net "out", 0 0, L_0x5c7c331528d0;  alias, 1 drivers
S_0x5c7c33033fb0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33033890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33034720_0 .net "in_a", 0 0, L_0x5c7c331528d0;  alias, 1 drivers
v0x5c7c330347c0_0 .net "out", 0 0, L_0x5c7c33152980;  alias, 1 drivers
S_0x5c7c330341d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33033fb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152980 .functor NAND 1, L_0x5c7c331528d0, L_0x5c7c331528d0, C4<1>, C4<1>;
v0x5c7c33034440_0 .net "in_a", 0 0, L_0x5c7c331528d0;  alias, 1 drivers
v0x5c7c33034530_0 .net "in_b", 0 0, L_0x5c7c331528d0;  alias, 1 drivers
v0x5c7c33034620_0 .net "out", 0 0, L_0x5c7c33152980;  alias, 1 drivers
S_0x5c7c33034ce0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33030d90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33035410_0 .net "in_a", 0 0, L_0x5c7c33152340;  alias, 1 drivers
v0x5c7c330354b0_0 .net "out", 0 0, L_0x5c7c331523f0;  alias, 1 drivers
S_0x5c7c33034eb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33034ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331523f0 .functor NAND 1, L_0x5c7c33152340, L_0x5c7c33152340, C4<1>, C4<1>;
v0x5c7c33035120_0 .net "in_a", 0 0, L_0x5c7c33152340;  alias, 1 drivers
v0x5c7c330351e0_0 .net "in_b", 0 0, L_0x5c7c33152340;  alias, 1 drivers
v0x5c7c33035330_0 .net "out", 0 0, L_0x5c7c331523f0;  alias, 1 drivers
S_0x5c7c330355b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33030d90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33035d80_0 .net "in_a", 0 0, L_0x5c7c33152660;  alias, 1 drivers
v0x5c7c33035e20_0 .net "out", 0 0, L_0x5c7c33152710;  alias, 1 drivers
S_0x5c7c33035820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330355b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152710 .functor NAND 1, L_0x5c7c33152660, L_0x5c7c33152660, C4<1>, C4<1>;
v0x5c7c33035a90_0 .net "in_a", 0 0, L_0x5c7c33152660;  alias, 1 drivers
v0x5c7c33035b50_0 .net "in_b", 0 0, L_0x5c7c33152660;  alias, 1 drivers
v0x5c7c33035ca0_0 .net "out", 0 0, L_0x5c7c33152710;  alias, 1 drivers
S_0x5c7c33035f20 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33030d90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330366c0_0 .net "in_a", 0 0, L_0x5c7c33152980;  alias, 1 drivers
v0x5c7c33036760_0 .net "out", 0 0, L_0x5c7c33152a30;  alias, 1 drivers
S_0x5c7c33036140 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33035f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33152a30 .functor NAND 1, L_0x5c7c33152980, L_0x5c7c33152980, C4<1>, C4<1>;
v0x5c7c330363b0_0 .net "in_a", 0 0, L_0x5c7c33152980;  alias, 1 drivers
v0x5c7c33036470_0 .net "in_b", 0 0, L_0x5c7c33152980;  alias, 1 drivers
v0x5c7c330365c0_0 .net "out", 0 0, L_0x5c7c33152a30;  alias, 1 drivers
S_0x5c7c33037700 .scope module, "mux_gate7" "Mux" 15 14, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33040a60_0 .net "in_a", 0 0, L_0x5c7c33153c30;  1 drivers
v0x5c7c33040b00_0 .net "in_b", 0 0, L_0x5c7c33153cd0;  1 drivers
v0x5c7c33040c10_0 .net "out", 0 0, L_0x5c7c33153a70;  1 drivers
v0x5c7c33040cb0_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33040d50_0 .net "sel_out", 0 0, L_0x5c7c33151eb0;  1 drivers
v0x5c7c33040ed0_0 .net "temp_a_out", 0 0, L_0x5c7c331530c0;  1 drivers
v0x5c7c33041080_0 .net "temp_b_out", 0 0, L_0x5c7c33153220;  1 drivers
S_0x5c7c33037900 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33037700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33038960_0 .net "in_a", 0 0, L_0x5c7c33153c30;  alias, 1 drivers
v0x5c7c33038a30_0 .net "in_b", 0 0, L_0x5c7c33151eb0;  alias, 1 drivers
v0x5c7c33038b00_0 .net "out", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
v0x5c7c33038c20_0 .net "temp_out", 0 0, L_0x5c7c33153010;  1 drivers
S_0x5c7c33037b70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33037900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153010 .functor NAND 1, L_0x5c7c33153c30, L_0x5c7c33151eb0, C4<1>, C4<1>;
v0x5c7c33037de0_0 .net "in_a", 0 0, L_0x5c7c33153c30;  alias, 1 drivers
v0x5c7c33037ec0_0 .net "in_b", 0 0, L_0x5c7c33151eb0;  alias, 1 drivers
v0x5c7c33037f80_0 .net "out", 0 0, L_0x5c7c33153010;  alias, 1 drivers
S_0x5c7c330380a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33037900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330387e0_0 .net "in_a", 0 0, L_0x5c7c33153010;  alias, 1 drivers
v0x5c7c33038880_0 .net "out", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
S_0x5c7c330382c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330380a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331530c0 .functor NAND 1, L_0x5c7c33153010, L_0x5c7c33153010, C4<1>, C4<1>;
v0x5c7c33038530_0 .net "in_a", 0 0, L_0x5c7c33153010;  alias, 1 drivers
v0x5c7c330385f0_0 .net "in_b", 0 0, L_0x5c7c33153010;  alias, 1 drivers
v0x5c7c330386e0_0 .net "out", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
S_0x5c7c33038ce0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33037700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33039cf0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33039d90_0 .net "in_b", 0 0, L_0x5c7c33153cd0;  alias, 1 drivers
v0x5c7c33039e80_0 .net "out", 0 0, L_0x5c7c33153220;  alias, 1 drivers
v0x5c7c33039fa0_0 .net "temp_out", 0 0, L_0x5c7c33153170;  1 drivers
S_0x5c7c33038ec0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33038ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153170 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33153cd0, C4<1>, C4<1>;
v0x5c7c33039130_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330391f0_0 .net "in_b", 0 0, L_0x5c7c33153cd0;  alias, 1 drivers
v0x5c7c330392b0_0 .net "out", 0 0, L_0x5c7c33153170;  alias, 1 drivers
S_0x5c7c330393d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33038ce0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33039b40_0 .net "in_a", 0 0, L_0x5c7c33153170;  alias, 1 drivers
v0x5c7c33039be0_0 .net "out", 0 0, L_0x5c7c33153220;  alias, 1 drivers
S_0x5c7c330395f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330393d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153220 .functor NAND 1, L_0x5c7c33153170, L_0x5c7c33153170, C4<1>, C4<1>;
v0x5c7c33039860_0 .net "in_a", 0 0, L_0x5c7c33153170;  alias, 1 drivers
v0x5c7c33039950_0 .net "in_b", 0 0, L_0x5c7c33153170;  alias, 1 drivers
v0x5c7c33039a40_0 .net "out", 0 0, L_0x5c7c33153220;  alias, 1 drivers
S_0x5c7c3303a060 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33037700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3303a760_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3303a800_0 .net "out", 0 0, L_0x5c7c33151eb0;  alias, 1 drivers
S_0x5c7c3303a230 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303a060;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33151eb0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c3303a480_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3303a540_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3303a600_0 .net "out", 0 0, L_0x5c7c33151eb0;  alias, 1 drivers
S_0x5c7c3303a900 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33037700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330403b0_0 .net "branch1_out", 0 0, L_0x5c7c33153430;  1 drivers
v0x5c7c330404e0_0 .net "branch2_out", 0 0, L_0x5c7c33153750;  1 drivers
v0x5c7c33040630_0 .net "in_a", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
v0x5c7c33040700_0 .net "in_b", 0 0, L_0x5c7c33153220;  alias, 1 drivers
v0x5c7c330407a0_0 .net "out", 0 0, L_0x5c7c33153a70;  alias, 1 drivers
v0x5c7c33040840_0 .net "temp1_out", 0 0, L_0x5c7c33153380;  1 drivers
v0x5c7c330408e0_0 .net "temp2_out", 0 0, L_0x5c7c331536a0;  1 drivers
v0x5c7c33040980_0 .net "temp3_out", 0 0, L_0x5c7c331539c0;  1 drivers
S_0x5c7c3303ab30 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c3303a900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3303bbf0_0 .net "in_a", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
v0x5c7c3303bc90_0 .net "in_b", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
v0x5c7c3303bd50_0 .net "out", 0 0, L_0x5c7c33153380;  alias, 1 drivers
v0x5c7c3303be70_0 .net "temp_out", 0 0, L_0x5c7c331532d0;  1 drivers
S_0x5c7c3303ada0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3303ab30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331532d0 .functor NAND 1, L_0x5c7c331530c0, L_0x5c7c331530c0, C4<1>, C4<1>;
v0x5c7c3303b010_0 .net "in_a", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
v0x5c7c3303b0d0_0 .net "in_b", 0 0, L_0x5c7c331530c0;  alias, 1 drivers
v0x5c7c3303b220_0 .net "out", 0 0, L_0x5c7c331532d0;  alias, 1 drivers
S_0x5c7c3303b320 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3303ab30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3303ba40_0 .net "in_a", 0 0, L_0x5c7c331532d0;  alias, 1 drivers
v0x5c7c3303bae0_0 .net "out", 0 0, L_0x5c7c33153380;  alias, 1 drivers
S_0x5c7c3303b4f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303b320;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153380 .functor NAND 1, L_0x5c7c331532d0, L_0x5c7c331532d0, C4<1>, C4<1>;
v0x5c7c3303b760_0 .net "in_a", 0 0, L_0x5c7c331532d0;  alias, 1 drivers
v0x5c7c3303b850_0 .net "in_b", 0 0, L_0x5c7c331532d0;  alias, 1 drivers
v0x5c7c3303b940_0 .net "out", 0 0, L_0x5c7c33153380;  alias, 1 drivers
S_0x5c7c3303bfe0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c3303a900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3303d010_0 .net "in_a", 0 0, L_0x5c7c33153220;  alias, 1 drivers
v0x5c7c3303d0b0_0 .net "in_b", 0 0, L_0x5c7c33153220;  alias, 1 drivers
v0x5c7c3303d170_0 .net "out", 0 0, L_0x5c7c331536a0;  alias, 1 drivers
v0x5c7c3303d290_0 .net "temp_out", 0 0, L_0x5c7c331535f0;  1 drivers
S_0x5c7c3303c1c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3303bfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331535f0 .functor NAND 1, L_0x5c7c33153220, L_0x5c7c33153220, C4<1>, C4<1>;
v0x5c7c3303c430_0 .net "in_a", 0 0, L_0x5c7c33153220;  alias, 1 drivers
v0x5c7c3303c4f0_0 .net "in_b", 0 0, L_0x5c7c33153220;  alias, 1 drivers
v0x5c7c3303c640_0 .net "out", 0 0, L_0x5c7c331535f0;  alias, 1 drivers
S_0x5c7c3303c740 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3303bfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3303ce60_0 .net "in_a", 0 0, L_0x5c7c331535f0;  alias, 1 drivers
v0x5c7c3303cf00_0 .net "out", 0 0, L_0x5c7c331536a0;  alias, 1 drivers
S_0x5c7c3303c910 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303c740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331536a0 .functor NAND 1, L_0x5c7c331535f0, L_0x5c7c331535f0, C4<1>, C4<1>;
v0x5c7c3303cb80_0 .net "in_a", 0 0, L_0x5c7c331535f0;  alias, 1 drivers
v0x5c7c3303cc70_0 .net "in_b", 0 0, L_0x5c7c331535f0;  alias, 1 drivers
v0x5c7c3303cd60_0 .net "out", 0 0, L_0x5c7c331536a0;  alias, 1 drivers
S_0x5c7c3303d400 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c3303a900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3303e440_0 .net "in_a", 0 0, L_0x5c7c33153430;  alias, 1 drivers
v0x5c7c3303e510_0 .net "in_b", 0 0, L_0x5c7c33153750;  alias, 1 drivers
v0x5c7c3303e5e0_0 .net "out", 0 0, L_0x5c7c331539c0;  alias, 1 drivers
v0x5c7c3303e700_0 .net "temp_out", 0 0, L_0x5c7c33153910;  1 drivers
S_0x5c7c3303d5e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3303d400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153910 .functor NAND 1, L_0x5c7c33153430, L_0x5c7c33153750, C4<1>, C4<1>;
v0x5c7c3303d830_0 .net "in_a", 0 0, L_0x5c7c33153430;  alias, 1 drivers
v0x5c7c3303d910_0 .net "in_b", 0 0, L_0x5c7c33153750;  alias, 1 drivers
v0x5c7c3303d9d0_0 .net "out", 0 0, L_0x5c7c33153910;  alias, 1 drivers
S_0x5c7c3303db20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3303d400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3303e290_0 .net "in_a", 0 0, L_0x5c7c33153910;  alias, 1 drivers
v0x5c7c3303e330_0 .net "out", 0 0, L_0x5c7c331539c0;  alias, 1 drivers
S_0x5c7c3303dd40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303db20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331539c0 .functor NAND 1, L_0x5c7c33153910, L_0x5c7c33153910, C4<1>, C4<1>;
v0x5c7c3303dfb0_0 .net "in_a", 0 0, L_0x5c7c33153910;  alias, 1 drivers
v0x5c7c3303e0a0_0 .net "in_b", 0 0, L_0x5c7c33153910;  alias, 1 drivers
v0x5c7c3303e190_0 .net "out", 0 0, L_0x5c7c331539c0;  alias, 1 drivers
S_0x5c7c3303e850 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c3303a900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3303ef80_0 .net "in_a", 0 0, L_0x5c7c33153380;  alias, 1 drivers
v0x5c7c3303f020_0 .net "out", 0 0, L_0x5c7c33153430;  alias, 1 drivers
S_0x5c7c3303ea20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303e850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153430 .functor NAND 1, L_0x5c7c33153380, L_0x5c7c33153380, C4<1>, C4<1>;
v0x5c7c3303ec90_0 .net "in_a", 0 0, L_0x5c7c33153380;  alias, 1 drivers
v0x5c7c3303ed50_0 .net "in_b", 0 0, L_0x5c7c33153380;  alias, 1 drivers
v0x5c7c3303eea0_0 .net "out", 0 0, L_0x5c7c33153430;  alias, 1 drivers
S_0x5c7c3303f120 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c3303a900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3303f8f0_0 .net "in_a", 0 0, L_0x5c7c331536a0;  alias, 1 drivers
v0x5c7c3303f990_0 .net "out", 0 0, L_0x5c7c33153750;  alias, 1 drivers
S_0x5c7c3303f390 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303f120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153750 .functor NAND 1, L_0x5c7c331536a0, L_0x5c7c331536a0, C4<1>, C4<1>;
v0x5c7c3303f600_0 .net "in_a", 0 0, L_0x5c7c331536a0;  alias, 1 drivers
v0x5c7c3303f6c0_0 .net "in_b", 0 0, L_0x5c7c331536a0;  alias, 1 drivers
v0x5c7c3303f810_0 .net "out", 0 0, L_0x5c7c33153750;  alias, 1 drivers
S_0x5c7c3303fa90 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c3303a900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33040230_0 .net "in_a", 0 0, L_0x5c7c331539c0;  alias, 1 drivers
v0x5c7c330402d0_0 .net "out", 0 0, L_0x5c7c33153a70;  alias, 1 drivers
S_0x5c7c3303fcb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3303fa90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153a70 .functor NAND 1, L_0x5c7c331539c0, L_0x5c7c331539c0, C4<1>, C4<1>;
v0x5c7c3303ff20_0 .net "in_a", 0 0, L_0x5c7c331539c0;  alias, 1 drivers
v0x5c7c3303ffe0_0 .net "in_b", 0 0, L_0x5c7c331539c0;  alias, 1 drivers
v0x5c7c33040130_0 .net "out", 0 0, L_0x5c7c33153a70;  alias, 1 drivers
S_0x5c7c33041270 .scope module, "mux_gate8" "Mux" 15 15, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c3304a5d0_0 .net "in_a", 0 0, L_0x5c7c33154ad0;  1 drivers
v0x5c7c3304a670_0 .net "in_b", 0 0, L_0x5c7c33154b70;  1 drivers
v0x5c7c3304a780_0 .net "out", 0 0, L_0x5c7c33154910;  1 drivers
v0x5c7c3304a820_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3304a8c0_0 .net "sel_out", 0 0, L_0x5c7c33153e00;  1 drivers
v0x5c7c3304aa40_0 .net "temp_a_out", 0 0, L_0x5c7c33153f60;  1 drivers
v0x5c7c3304abf0_0 .net "temp_b_out", 0 0, L_0x5c7c331540c0;  1 drivers
S_0x5c7c33041470 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33041270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330424d0_0 .net "in_a", 0 0, L_0x5c7c33154ad0;  alias, 1 drivers
v0x5c7c330425a0_0 .net "in_b", 0 0, L_0x5c7c33153e00;  alias, 1 drivers
v0x5c7c33042670_0 .net "out", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
v0x5c7c33042790_0 .net "temp_out", 0 0, L_0x5c7c33153eb0;  1 drivers
S_0x5c7c330416e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33041470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153eb0 .functor NAND 1, L_0x5c7c33154ad0, L_0x5c7c33153e00, C4<1>, C4<1>;
v0x5c7c33041950_0 .net "in_a", 0 0, L_0x5c7c33154ad0;  alias, 1 drivers
v0x5c7c33041a30_0 .net "in_b", 0 0, L_0x5c7c33153e00;  alias, 1 drivers
v0x5c7c33041af0_0 .net "out", 0 0, L_0x5c7c33153eb0;  alias, 1 drivers
S_0x5c7c33041c10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33041470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33042350_0 .net "in_a", 0 0, L_0x5c7c33153eb0;  alias, 1 drivers
v0x5c7c330423f0_0 .net "out", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
S_0x5c7c33041e30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33041c10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153f60 .functor NAND 1, L_0x5c7c33153eb0, L_0x5c7c33153eb0, C4<1>, C4<1>;
v0x5c7c330420a0_0 .net "in_a", 0 0, L_0x5c7c33153eb0;  alias, 1 drivers
v0x5c7c33042160_0 .net "in_b", 0 0, L_0x5c7c33153eb0;  alias, 1 drivers
v0x5c7c33042250_0 .net "out", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
S_0x5c7c33042850 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33041270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33043860_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33043900_0 .net "in_b", 0 0, L_0x5c7c33154b70;  alias, 1 drivers
v0x5c7c330439f0_0 .net "out", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
v0x5c7c33043b10_0 .net "temp_out", 0 0, L_0x5c7c33154010;  1 drivers
S_0x5c7c33042a30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33042850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154010 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33154b70, C4<1>, C4<1>;
v0x5c7c33042ca0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33042d60_0 .net "in_b", 0 0, L_0x5c7c33154b70;  alias, 1 drivers
v0x5c7c33042e20_0 .net "out", 0 0, L_0x5c7c33154010;  alias, 1 drivers
S_0x5c7c33042f40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33042850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330436b0_0 .net "in_a", 0 0, L_0x5c7c33154010;  alias, 1 drivers
v0x5c7c33043750_0 .net "out", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
S_0x5c7c33043160 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33042f40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331540c0 .functor NAND 1, L_0x5c7c33154010, L_0x5c7c33154010, C4<1>, C4<1>;
v0x5c7c330433d0_0 .net "in_a", 0 0, L_0x5c7c33154010;  alias, 1 drivers
v0x5c7c330434c0_0 .net "in_b", 0 0, L_0x5c7c33154010;  alias, 1 drivers
v0x5c7c330435b0_0 .net "out", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
S_0x5c7c33043bd0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33041270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330442d0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33044370_0 .net "out", 0 0, L_0x5c7c33153e00;  alias, 1 drivers
S_0x5c7c33043da0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33043bd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33153e00 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c33043ff0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c330440b0_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33044170_0 .net "out", 0 0, L_0x5c7c33153e00;  alias, 1 drivers
S_0x5c7c33044470 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33041270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33049f20_0 .net "branch1_out", 0 0, L_0x5c7c331542d0;  1 drivers
v0x5c7c3304a050_0 .net "branch2_out", 0 0, L_0x5c7c331545f0;  1 drivers
v0x5c7c3304a1a0_0 .net "in_a", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
v0x5c7c3304a270_0 .net "in_b", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
v0x5c7c3304a310_0 .net "out", 0 0, L_0x5c7c33154910;  alias, 1 drivers
v0x5c7c3304a3b0_0 .net "temp1_out", 0 0, L_0x5c7c33154220;  1 drivers
v0x5c7c3304a450_0 .net "temp2_out", 0 0, L_0x5c7c33154540;  1 drivers
v0x5c7c3304a4f0_0 .net "temp3_out", 0 0, L_0x5c7c33154860;  1 drivers
S_0x5c7c330446a0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33044470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33045760_0 .net "in_a", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
v0x5c7c33045800_0 .net "in_b", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
v0x5c7c330458c0_0 .net "out", 0 0, L_0x5c7c33154220;  alias, 1 drivers
v0x5c7c330459e0_0 .net "temp_out", 0 0, L_0x5c7c33154170;  1 drivers
S_0x5c7c33044910 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330446a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154170 .functor NAND 1, L_0x5c7c33153f60, L_0x5c7c33153f60, C4<1>, C4<1>;
v0x5c7c33044b80_0 .net "in_a", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
v0x5c7c33044c40_0 .net "in_b", 0 0, L_0x5c7c33153f60;  alias, 1 drivers
v0x5c7c33044d90_0 .net "out", 0 0, L_0x5c7c33154170;  alias, 1 drivers
S_0x5c7c33044e90 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330446a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330455b0_0 .net "in_a", 0 0, L_0x5c7c33154170;  alias, 1 drivers
v0x5c7c33045650_0 .net "out", 0 0, L_0x5c7c33154220;  alias, 1 drivers
S_0x5c7c33045060 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33044e90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154220 .functor NAND 1, L_0x5c7c33154170, L_0x5c7c33154170, C4<1>, C4<1>;
v0x5c7c330452d0_0 .net "in_a", 0 0, L_0x5c7c33154170;  alias, 1 drivers
v0x5c7c330453c0_0 .net "in_b", 0 0, L_0x5c7c33154170;  alias, 1 drivers
v0x5c7c330454b0_0 .net "out", 0 0, L_0x5c7c33154220;  alias, 1 drivers
S_0x5c7c33045b50 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33044470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33046b80_0 .net "in_a", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
v0x5c7c33046c20_0 .net "in_b", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
v0x5c7c33046ce0_0 .net "out", 0 0, L_0x5c7c33154540;  alias, 1 drivers
v0x5c7c33046e00_0 .net "temp_out", 0 0, L_0x5c7c33154490;  1 drivers
S_0x5c7c33045d30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33045b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154490 .functor NAND 1, L_0x5c7c331540c0, L_0x5c7c331540c0, C4<1>, C4<1>;
v0x5c7c33045fa0_0 .net "in_a", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
v0x5c7c33046060_0 .net "in_b", 0 0, L_0x5c7c331540c0;  alias, 1 drivers
v0x5c7c330461b0_0 .net "out", 0 0, L_0x5c7c33154490;  alias, 1 drivers
S_0x5c7c330462b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33045b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330469d0_0 .net "in_a", 0 0, L_0x5c7c33154490;  alias, 1 drivers
v0x5c7c33046a70_0 .net "out", 0 0, L_0x5c7c33154540;  alias, 1 drivers
S_0x5c7c33046480 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330462b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154540 .functor NAND 1, L_0x5c7c33154490, L_0x5c7c33154490, C4<1>, C4<1>;
v0x5c7c330466f0_0 .net "in_a", 0 0, L_0x5c7c33154490;  alias, 1 drivers
v0x5c7c330467e0_0 .net "in_b", 0 0, L_0x5c7c33154490;  alias, 1 drivers
v0x5c7c330468d0_0 .net "out", 0 0, L_0x5c7c33154540;  alias, 1 drivers
S_0x5c7c33046f70 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33044470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33047fb0_0 .net "in_a", 0 0, L_0x5c7c331542d0;  alias, 1 drivers
v0x5c7c33048080_0 .net "in_b", 0 0, L_0x5c7c331545f0;  alias, 1 drivers
v0x5c7c33048150_0 .net "out", 0 0, L_0x5c7c33154860;  alias, 1 drivers
v0x5c7c33048270_0 .net "temp_out", 0 0, L_0x5c7c331547b0;  1 drivers
S_0x5c7c33047150 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33046f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331547b0 .functor NAND 1, L_0x5c7c331542d0, L_0x5c7c331545f0, C4<1>, C4<1>;
v0x5c7c330473a0_0 .net "in_a", 0 0, L_0x5c7c331542d0;  alias, 1 drivers
v0x5c7c33047480_0 .net "in_b", 0 0, L_0x5c7c331545f0;  alias, 1 drivers
v0x5c7c33047540_0 .net "out", 0 0, L_0x5c7c331547b0;  alias, 1 drivers
S_0x5c7c33047690 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33046f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33047e00_0 .net "in_a", 0 0, L_0x5c7c331547b0;  alias, 1 drivers
v0x5c7c33047ea0_0 .net "out", 0 0, L_0x5c7c33154860;  alias, 1 drivers
S_0x5c7c330478b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33047690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154860 .functor NAND 1, L_0x5c7c331547b0, L_0x5c7c331547b0, C4<1>, C4<1>;
v0x5c7c33047b20_0 .net "in_a", 0 0, L_0x5c7c331547b0;  alias, 1 drivers
v0x5c7c33047c10_0 .net "in_b", 0 0, L_0x5c7c331547b0;  alias, 1 drivers
v0x5c7c33047d00_0 .net "out", 0 0, L_0x5c7c33154860;  alias, 1 drivers
S_0x5c7c330483c0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33044470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33048af0_0 .net "in_a", 0 0, L_0x5c7c33154220;  alias, 1 drivers
v0x5c7c33048b90_0 .net "out", 0 0, L_0x5c7c331542d0;  alias, 1 drivers
S_0x5c7c33048590 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330483c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331542d0 .functor NAND 1, L_0x5c7c33154220, L_0x5c7c33154220, C4<1>, C4<1>;
v0x5c7c33048800_0 .net "in_a", 0 0, L_0x5c7c33154220;  alias, 1 drivers
v0x5c7c330488c0_0 .net "in_b", 0 0, L_0x5c7c33154220;  alias, 1 drivers
v0x5c7c33048a10_0 .net "out", 0 0, L_0x5c7c331542d0;  alias, 1 drivers
S_0x5c7c33048c90 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33044470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33049460_0 .net "in_a", 0 0, L_0x5c7c33154540;  alias, 1 drivers
v0x5c7c33049500_0 .net "out", 0 0, L_0x5c7c331545f0;  alias, 1 drivers
S_0x5c7c33048f00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33048c90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331545f0 .functor NAND 1, L_0x5c7c33154540, L_0x5c7c33154540, C4<1>, C4<1>;
v0x5c7c33049170_0 .net "in_a", 0 0, L_0x5c7c33154540;  alias, 1 drivers
v0x5c7c33049230_0 .net "in_b", 0 0, L_0x5c7c33154540;  alias, 1 drivers
v0x5c7c33049380_0 .net "out", 0 0, L_0x5c7c331545f0;  alias, 1 drivers
S_0x5c7c33049600 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33044470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33049da0_0 .net "in_a", 0 0, L_0x5c7c33154860;  alias, 1 drivers
v0x5c7c33049e40_0 .net "out", 0 0, L_0x5c7c33154910;  alias, 1 drivers
S_0x5c7c33049820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33049600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154910 .functor NAND 1, L_0x5c7c33154860, L_0x5c7c33154860, C4<1>, C4<1>;
v0x5c7c33049a90_0 .net "in_a", 0 0, L_0x5c7c33154860;  alias, 1 drivers
v0x5c7c33049b50_0 .net "in_b", 0 0, L_0x5c7c33154860;  alias, 1 drivers
v0x5c7c33049ca0_0 .net "out", 0 0, L_0x5c7c33154910;  alias, 1 drivers
S_0x5c7c3304ade0 .scope module, "mux_gate9" "Mux" 15 16, 16 3 0, S_0x5c7c32fb86e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33054140_0 .net "in_a", 0 0, L_0x5c7c33155980;  1 drivers
v0x5c7c330541e0_0 .net "in_b", 0 0, L_0x5c7c33155a20;  1 drivers
v0x5c7c330542f0_0 .net "out", 0 0, L_0x5c7c331557c0;  1 drivers
v0x5c7c33054390_0 .net "sel", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c33054430_0 .net "sel_out", 0 0, L_0x5c7c33154cb0;  1 drivers
v0x5c7c330545b0_0 .net "temp_a_out", 0 0, L_0x5c7c33154e10;  1 drivers
v0x5c7c33054760_0 .net "temp_b_out", 0 0, L_0x5c7c33154f70;  1 drivers
S_0x5c7c3304afe0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c3304ade0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3304c040_0 .net "in_a", 0 0, L_0x5c7c33155980;  alias, 1 drivers
v0x5c7c3304c110_0 .net "in_b", 0 0, L_0x5c7c33154cb0;  alias, 1 drivers
v0x5c7c3304c1e0_0 .net "out", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
v0x5c7c3304c300_0 .net "temp_out", 0 0, L_0x5c7c33154d60;  1 drivers
S_0x5c7c3304b250 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3304afe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154d60 .functor NAND 1, L_0x5c7c33155980, L_0x5c7c33154cb0, C4<1>, C4<1>;
v0x5c7c3304b4c0_0 .net "in_a", 0 0, L_0x5c7c33155980;  alias, 1 drivers
v0x5c7c3304b5a0_0 .net "in_b", 0 0, L_0x5c7c33154cb0;  alias, 1 drivers
v0x5c7c3304b660_0 .net "out", 0 0, L_0x5c7c33154d60;  alias, 1 drivers
S_0x5c7c3304b780 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3304afe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3304bec0_0 .net "in_a", 0 0, L_0x5c7c33154d60;  alias, 1 drivers
v0x5c7c3304bf60_0 .net "out", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
S_0x5c7c3304b9a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3304b780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154e10 .functor NAND 1, L_0x5c7c33154d60, L_0x5c7c33154d60, C4<1>, C4<1>;
v0x5c7c3304bc10_0 .net "in_a", 0 0, L_0x5c7c33154d60;  alias, 1 drivers
v0x5c7c3304bcd0_0 .net "in_b", 0 0, L_0x5c7c33154d60;  alias, 1 drivers
v0x5c7c3304bdc0_0 .net "out", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
S_0x5c7c3304c3c0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c3304ade0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3304d3d0_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3304d470_0 .net "in_b", 0 0, L_0x5c7c33155a20;  alias, 1 drivers
v0x5c7c3304d560_0 .net "out", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
v0x5c7c3304d680_0 .net "temp_out", 0 0, L_0x5c7c33154ec0;  1 drivers
S_0x5c7c3304c5a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3304c3c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154ec0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c33155a20, C4<1>, C4<1>;
v0x5c7c3304c810_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3304c8d0_0 .net "in_b", 0 0, L_0x5c7c33155a20;  alias, 1 drivers
v0x5c7c3304c990_0 .net "out", 0 0, L_0x5c7c33154ec0;  alias, 1 drivers
S_0x5c7c3304cab0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3304c3c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3304d220_0 .net "in_a", 0 0, L_0x5c7c33154ec0;  alias, 1 drivers
v0x5c7c3304d2c0_0 .net "out", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
S_0x5c7c3304ccd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3304cab0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154f70 .functor NAND 1, L_0x5c7c33154ec0, L_0x5c7c33154ec0, C4<1>, C4<1>;
v0x5c7c3304cf40_0 .net "in_a", 0 0, L_0x5c7c33154ec0;  alias, 1 drivers
v0x5c7c3304d030_0 .net "in_b", 0 0, L_0x5c7c33154ec0;  alias, 1 drivers
v0x5c7c3304d120_0 .net "out", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
S_0x5c7c3304d740 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c3304ade0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3304de40_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3304dee0_0 .net "out", 0 0, L_0x5c7c33154cb0;  alias, 1 drivers
S_0x5c7c3304d910 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3304d740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33154cb0 .functor NAND 1, L_0x5c7c3315b570, L_0x5c7c3315b570, C4<1>, C4<1>;
v0x5c7c3304db60_0 .net "in_a", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3304dc20_0 .net "in_b", 0 0, L_0x5c7c3315b570;  alias, 1 drivers
v0x5c7c3304dce0_0 .net "out", 0 0, L_0x5c7c33154cb0;  alias, 1 drivers
S_0x5c7c3304dfe0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c3304ade0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33053a90_0 .net "branch1_out", 0 0, L_0x5c7c33155180;  1 drivers
v0x5c7c33053bc0_0 .net "branch2_out", 0 0, L_0x5c7c331554a0;  1 drivers
v0x5c7c33053d10_0 .net "in_a", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
v0x5c7c33053de0_0 .net "in_b", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
v0x5c7c33053e80_0 .net "out", 0 0, L_0x5c7c331557c0;  alias, 1 drivers
v0x5c7c33053f20_0 .net "temp1_out", 0 0, L_0x5c7c331550d0;  1 drivers
v0x5c7c33053fc0_0 .net "temp2_out", 0 0, L_0x5c7c331553f0;  1 drivers
v0x5c7c33054060_0 .net "temp3_out", 0 0, L_0x5c7c33155710;  1 drivers
S_0x5c7c3304e210 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c3304dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3304f2d0_0 .net "in_a", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
v0x5c7c3304f370_0 .net "in_b", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
v0x5c7c3304f430_0 .net "out", 0 0, L_0x5c7c331550d0;  alias, 1 drivers
v0x5c7c3304f550_0 .net "temp_out", 0 0, L_0x5c7c33155020;  1 drivers
S_0x5c7c3304e480 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3304e210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33155020 .functor NAND 1, L_0x5c7c33154e10, L_0x5c7c33154e10, C4<1>, C4<1>;
v0x5c7c3304e6f0_0 .net "in_a", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
v0x5c7c3304e7b0_0 .net "in_b", 0 0, L_0x5c7c33154e10;  alias, 1 drivers
v0x5c7c3304e900_0 .net "out", 0 0, L_0x5c7c33155020;  alias, 1 drivers
S_0x5c7c3304ea00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3304e210;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3304f120_0 .net "in_a", 0 0, L_0x5c7c33155020;  alias, 1 drivers
v0x5c7c3304f1c0_0 .net "out", 0 0, L_0x5c7c331550d0;  alias, 1 drivers
S_0x5c7c3304ebd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3304ea00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331550d0 .functor NAND 1, L_0x5c7c33155020, L_0x5c7c33155020, C4<1>, C4<1>;
v0x5c7c3304ee40_0 .net "in_a", 0 0, L_0x5c7c33155020;  alias, 1 drivers
v0x5c7c3304ef30_0 .net "in_b", 0 0, L_0x5c7c33155020;  alias, 1 drivers
v0x5c7c3304f020_0 .net "out", 0 0, L_0x5c7c331550d0;  alias, 1 drivers
S_0x5c7c3304f6c0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c3304dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330506f0_0 .net "in_a", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
v0x5c7c33050790_0 .net "in_b", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
v0x5c7c33050850_0 .net "out", 0 0, L_0x5c7c331553f0;  alias, 1 drivers
v0x5c7c33050970_0 .net "temp_out", 0 0, L_0x5c7c33155340;  1 drivers
S_0x5c7c3304f8a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3304f6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33155340 .functor NAND 1, L_0x5c7c33154f70, L_0x5c7c33154f70, C4<1>, C4<1>;
v0x5c7c3304fb10_0 .net "in_a", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
v0x5c7c3304fbd0_0 .net "in_b", 0 0, L_0x5c7c33154f70;  alias, 1 drivers
v0x5c7c3304fd20_0 .net "out", 0 0, L_0x5c7c33155340;  alias, 1 drivers
S_0x5c7c3304fe20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3304f6c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33050540_0 .net "in_a", 0 0, L_0x5c7c33155340;  alias, 1 drivers
v0x5c7c330505e0_0 .net "out", 0 0, L_0x5c7c331553f0;  alias, 1 drivers
S_0x5c7c3304fff0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3304fe20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331553f0 .functor NAND 1, L_0x5c7c33155340, L_0x5c7c33155340, C4<1>, C4<1>;
v0x5c7c33050260_0 .net "in_a", 0 0, L_0x5c7c33155340;  alias, 1 drivers
v0x5c7c33050350_0 .net "in_b", 0 0, L_0x5c7c33155340;  alias, 1 drivers
v0x5c7c33050440_0 .net "out", 0 0, L_0x5c7c331553f0;  alias, 1 drivers
S_0x5c7c33050ae0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c3304dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33051b20_0 .net "in_a", 0 0, L_0x5c7c33155180;  alias, 1 drivers
v0x5c7c33051bf0_0 .net "in_b", 0 0, L_0x5c7c331554a0;  alias, 1 drivers
v0x5c7c33051cc0_0 .net "out", 0 0, L_0x5c7c33155710;  alias, 1 drivers
v0x5c7c33051de0_0 .net "temp_out", 0 0, L_0x5c7c33155660;  1 drivers
S_0x5c7c33050cc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33050ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33155660 .functor NAND 1, L_0x5c7c33155180, L_0x5c7c331554a0, C4<1>, C4<1>;
v0x5c7c33050f10_0 .net "in_a", 0 0, L_0x5c7c33155180;  alias, 1 drivers
v0x5c7c33050ff0_0 .net "in_b", 0 0, L_0x5c7c331554a0;  alias, 1 drivers
v0x5c7c330510b0_0 .net "out", 0 0, L_0x5c7c33155660;  alias, 1 drivers
S_0x5c7c33051200 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33050ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33051970_0 .net "in_a", 0 0, L_0x5c7c33155660;  alias, 1 drivers
v0x5c7c33051a10_0 .net "out", 0 0, L_0x5c7c33155710;  alias, 1 drivers
S_0x5c7c33051420 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33051200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33155710 .functor NAND 1, L_0x5c7c33155660, L_0x5c7c33155660, C4<1>, C4<1>;
v0x5c7c33051690_0 .net "in_a", 0 0, L_0x5c7c33155660;  alias, 1 drivers
v0x5c7c33051780_0 .net "in_b", 0 0, L_0x5c7c33155660;  alias, 1 drivers
v0x5c7c33051870_0 .net "out", 0 0, L_0x5c7c33155710;  alias, 1 drivers
S_0x5c7c33051f30 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c3304dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33052660_0 .net "in_a", 0 0, L_0x5c7c331550d0;  alias, 1 drivers
v0x5c7c33052700_0 .net "out", 0 0, L_0x5c7c33155180;  alias, 1 drivers
S_0x5c7c33052100 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33051f30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33155180 .functor NAND 1, L_0x5c7c331550d0, L_0x5c7c331550d0, C4<1>, C4<1>;
v0x5c7c33052370_0 .net "in_a", 0 0, L_0x5c7c331550d0;  alias, 1 drivers
v0x5c7c33052430_0 .net "in_b", 0 0, L_0x5c7c331550d0;  alias, 1 drivers
v0x5c7c33052580_0 .net "out", 0 0, L_0x5c7c33155180;  alias, 1 drivers
S_0x5c7c33052800 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c3304dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33052fd0_0 .net "in_a", 0 0, L_0x5c7c331553f0;  alias, 1 drivers
v0x5c7c33053070_0 .net "out", 0 0, L_0x5c7c331554a0;  alias, 1 drivers
S_0x5c7c33052a70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33052800;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331554a0 .functor NAND 1, L_0x5c7c331553f0, L_0x5c7c331553f0, C4<1>, C4<1>;
v0x5c7c33052ce0_0 .net "in_a", 0 0, L_0x5c7c331553f0;  alias, 1 drivers
v0x5c7c33052da0_0 .net "in_b", 0 0, L_0x5c7c331553f0;  alias, 1 drivers
v0x5c7c33052ef0_0 .net "out", 0 0, L_0x5c7c331554a0;  alias, 1 drivers
S_0x5c7c33053170 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c3304dfe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33053910_0 .net "in_a", 0 0, L_0x5c7c33155710;  alias, 1 drivers
v0x5c7c330539b0_0 .net "out", 0 0, L_0x5c7c331557c0;  alias, 1 drivers
S_0x5c7c33053390 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33053170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331557c0 .functor NAND 1, L_0x5c7c33155710, L_0x5c7c33155710, C4<1>, C4<1>;
v0x5c7c33053600_0 .net "in_a", 0 0, L_0x5c7c33155710;  alias, 1 drivers
v0x5c7c330536c0_0 .net "in_b", 0 0, L_0x5c7c33155710;  alias, 1 drivers
v0x5c7c33053810_0 .net "out", 0 0, L_0x5c7c331557c0;  alias, 1 drivers
S_0x5c7c33054df0 .scope module, "mux16_gate3" "Mux16" 14 17, 15 3 0, S_0x5c7c32cac1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 16 "in_a";
    .port_info 1 /INPUT 16 "in_b";
    .port_info 2 /OUTPUT 16 "out";
    .port_info 3 /INPUT 1 "sel";
L_0x5c7c33169f80 .functor BUFZ 16, L_0x5c7c33169ee0, C4<0000000000000000>, C4<0000000000000000>, C4<0000000000000000>;
v0x5c7c33111070_0 .net "in_a", 15 0, L_0x5c7c3314c880;  alias, 1 drivers
v0x5c7c33111150_0 .net "in_b", 15 0, L_0x5c7c3315b4e0;  alias, 1 drivers
v0x5c7c331111f0_0 .net "out", 15 0, L_0x5c7c33169f80;  alias, 1 drivers
v0x5c7c33111290_0 .net "sel", 0 0, L_0x5c7c33169ff0;  1 drivers
v0x5c7c33111330_0 .net/s "tmp_out", 15 0, L_0x5c7c33169ee0;  1 drivers
L_0x5c7c3315c2e0 .part L_0x5c7c3314c880, 0, 1;
L_0x5c7c3315c3a0 .part L_0x5c7c3315b4e0, 0, 1;
L_0x5c7c3315d110 .part L_0x5c7c3314c880, 1, 1;
L_0x5c7c3315d1b0 .part L_0x5c7c3315b4e0, 1, 1;
L_0x5c7c3315df00 .part L_0x5c7c3314c880, 2, 1;
L_0x5c7c3315dfa0 .part L_0x5c7c3315b4e0, 2, 1;
L_0x5c7c3315ed50 .part L_0x5c7c3314c880, 3, 1;
L_0x5c7c3315edf0 .part L_0x5c7c3315b4e0, 3, 1;
L_0x5c7c3315fb60 .part L_0x5c7c3314c880, 4, 1;
L_0x5c7c3315fd10 .part L_0x5c7c3315b4e0, 4, 1;
L_0x5c7c33160bf0 .part L_0x5c7c3314c880, 5, 1;
L_0x5c7c33160c90 .part L_0x5c7c3315b4e0, 5, 1;
L_0x5c7c33161a70 .part L_0x5c7c3314c880, 6, 1;
L_0x5c7c33161b10 .part L_0x5c7c3315b4e0, 6, 1;
L_0x5c7c33162890 .part L_0x5c7c3314c880, 7, 1;
L_0x5c7c33162930 .part L_0x5c7c3315b4e0, 7, 1;
L_0x5c7c33163730 .part L_0x5c7c3314c880, 8, 1;
L_0x5c7c331637d0 .part L_0x5c7c3315b4e0, 8, 1;
L_0x5c7c331645e0 .part L_0x5c7c3314c880, 9, 1;
L_0x5c7c33164680 .part L_0x5c7c3315b4e0, 9, 1;
L_0x5c7c33163870 .part L_0x5c7c3314c880, 10, 1;
L_0x5c7c33165be0 .part L_0x5c7c3315b4e0, 10, 1;
L_0x5c7c33166690 .part L_0x5c7c3314c880, 11, 1;
L_0x5c7c33166730 .part L_0x5c7c3315b4e0, 11, 1;
L_0x5c7c331671f0 .part L_0x5c7c3314c880, 12, 1;
L_0x5c7c331674a0 .part L_0x5c7c3315b4e0, 12, 1;
L_0x5c7c33167f60 .part L_0x5c7c3314c880, 13, 1;
L_0x5c7c33168000 .part L_0x5c7c3315b4e0, 13, 1;
L_0x5c7c33168d80 .part L_0x5c7c3314c880, 14, 1;
L_0x5c7c33168e20 .part L_0x5c7c3315b4e0, 14, 1;
L_0x5c7c33169c90 .part L_0x5c7c3314c880, 15, 1;
L_0x5c7c33169d30 .part L_0x5c7c3315b4e0, 15, 1;
LS_0x5c7c33169ee0_0_0 .concat8 [ 1 1 1 1], L_0x5c7c3315c120, L_0x5c7c3315cf50, L_0x5c7c3315dd40, L_0x5c7c3315eb90;
LS_0x5c7c33169ee0_0_4 .concat8 [ 1 1 1 1], L_0x5c7c3315f9a0, L_0x5c7c33160a30, L_0x5c7c331618b0, L_0x5c7c331626d0;
LS_0x5c7c33169ee0_0_8 .concat8 [ 1 1 1 1], L_0x5c7c33163570, L_0x5c7c33164420, L_0x5c7c33165a60, L_0x5c7c33166510;
LS_0x5c7c33169ee0_0_12 .concat8 [ 1 1 1 1], L_0x5c7c33167070, L_0x5c7c33167de0, L_0x5c7c33168bc0, L_0x5c7c33169ad0;
L_0x5c7c33169ee0 .concat8 [ 4 4 4 4], LS_0x5c7c33169ee0_0_0, LS_0x5c7c33169ee0_0_4, LS_0x5c7c33169ee0_0_8, LS_0x5c7c33169ee0_0_12;
S_0x5c7c33055040 .scope module, "mux_gate0" "Mux" 15 7, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c3307e4e0_0 .net "in_a", 0 0, L_0x5c7c3315c2e0;  1 drivers
v0x5c7c3307e580_0 .net "in_b", 0 0, L_0x5c7c3315c3a0;  1 drivers
v0x5c7c3307e690_0 .net "out", 0 0, L_0x5c7c3315c120;  1 drivers
v0x5c7c3307e730_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3307e7d0_0 .net "sel_out", 0 0, L_0x5c7c3315b610;  1 drivers
v0x5c7c3307e950_0 .net "temp_a_out", 0 0, L_0x5c7c3315b770;  1 drivers
v0x5c7c3307eb00_0 .net "temp_b_out", 0 0, L_0x5c7c3315b8d0;  1 drivers
S_0x5c7c33055290 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33055040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33056350_0 .net "in_a", 0 0, L_0x5c7c3315c2e0;  alias, 1 drivers
v0x5c7c33056420_0 .net "in_b", 0 0, L_0x5c7c3315b610;  alias, 1 drivers
v0x5c7c330564f0_0 .net "out", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
v0x5c7c33056610_0 .net "temp_out", 0 0, L_0x5c7c3315b6c0;  1 drivers
S_0x5c7c33055500 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33055290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b6c0 .functor NAND 1, L_0x5c7c3315c2e0, L_0x5c7c3315b610, C4<1>, C4<1>;
v0x5c7c33055770_0 .net "in_a", 0 0, L_0x5c7c3315c2e0;  alias, 1 drivers
v0x5c7c33055850_0 .net "in_b", 0 0, L_0x5c7c3315b610;  alias, 1 drivers
v0x5c7c33055910_0 .net "out", 0 0, L_0x5c7c3315b6c0;  alias, 1 drivers
S_0x5c7c33055a30 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33055290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330561a0_0 .net "in_a", 0 0, L_0x5c7c3315b6c0;  alias, 1 drivers
v0x5c7c33056240_0 .net "out", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
S_0x5c7c33055c50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33055a30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b770 .functor NAND 1, L_0x5c7c3315b6c0, L_0x5c7c3315b6c0, C4<1>, C4<1>;
v0x5c7c33055ec0_0 .net "in_a", 0 0, L_0x5c7c3315b6c0;  alias, 1 drivers
v0x5c7c33055fb0_0 .net "in_b", 0 0, L_0x5c7c3315b6c0;  alias, 1 drivers
v0x5c7c330560a0_0 .net "out", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
S_0x5c7c330566d0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33055040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33057700_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330577d0_0 .net "in_b", 0 0, L_0x5c7c3315c3a0;  alias, 1 drivers
v0x5c7c330578a0_0 .net "out", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
v0x5c7c330579c0_0 .net "temp_out", 0 0, L_0x5c7c3315b820;  1 drivers
S_0x5c7c330568b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330566d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b820 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c3315c3a0, C4<1>, C4<1>;
v0x5c7c33056b20_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33056c00_0 .net "in_b", 0 0, L_0x5c7c3315c3a0;  alias, 1 drivers
v0x5c7c33056cc0_0 .net "out", 0 0, L_0x5c7c3315b820;  alias, 1 drivers
S_0x5c7c33056de0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330566d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33057550_0 .net "in_a", 0 0, L_0x5c7c3315b820;  alias, 1 drivers
v0x5c7c330575f0_0 .net "out", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
S_0x5c7c33057000 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33056de0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b8d0 .functor NAND 1, L_0x5c7c3315b820, L_0x5c7c3315b820, C4<1>, C4<1>;
v0x5c7c33057270_0 .net "in_a", 0 0, L_0x5c7c3315b820;  alias, 1 drivers
v0x5c7c33057360_0 .net "in_b", 0 0, L_0x5c7c3315b820;  alias, 1 drivers
v0x5c7c33057450_0 .net "out", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
S_0x5c7c33057a80 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33055040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330581a0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330582d0_0 .net "out", 0 0, L_0x5c7c3315b610;  alias, 1 drivers
S_0x5c7c33057c50 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33057a80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b610 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c33057ea0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33057fb0_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33058070_0 .net "out", 0 0, L_0x5c7c3315b610;  alias, 1 drivers
S_0x5c7c330583d0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33055040;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3307de30_0 .net "branch1_out", 0 0, L_0x5c7c3315bae0;  1 drivers
v0x5c7c3307df60_0 .net "branch2_out", 0 0, L_0x5c7c3315be00;  1 drivers
v0x5c7c3307e0b0_0 .net "in_a", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
v0x5c7c3307e180_0 .net "in_b", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
v0x5c7c3307e220_0 .net "out", 0 0, L_0x5c7c3315c120;  alias, 1 drivers
v0x5c7c3307e2c0_0 .net "temp1_out", 0 0, L_0x5c7c3315ba30;  1 drivers
v0x5c7c3307e360_0 .net "temp2_out", 0 0, L_0x5c7c3315bd50;  1 drivers
v0x5c7c3307e400_0 .net "temp3_out", 0 0, L_0x5c7c3315c070;  1 drivers
S_0x5c7c330585b0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330583d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33059670_0 .net "in_a", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
v0x5c7c33059710_0 .net "in_b", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
v0x5c7c330597d0_0 .net "out", 0 0, L_0x5c7c3315ba30;  alias, 1 drivers
v0x5c7c330598f0_0 .net "temp_out", 0 0, L_0x5c7c3315b980;  1 drivers
S_0x5c7c33058820 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330585b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315b980 .functor NAND 1, L_0x5c7c3315b770, L_0x5c7c3315b770, C4<1>, C4<1>;
v0x5c7c33058a90_0 .net "in_a", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
v0x5c7c33058b50_0 .net "in_b", 0 0, L_0x5c7c3315b770;  alias, 1 drivers
v0x5c7c33058ca0_0 .net "out", 0 0, L_0x5c7c3315b980;  alias, 1 drivers
S_0x5c7c33058da0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330585b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330594c0_0 .net "in_a", 0 0, L_0x5c7c3315b980;  alias, 1 drivers
v0x5c7c33059560_0 .net "out", 0 0, L_0x5c7c3315ba30;  alias, 1 drivers
S_0x5c7c33058f70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33058da0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ba30 .functor NAND 1, L_0x5c7c3315b980, L_0x5c7c3315b980, C4<1>, C4<1>;
v0x5c7c330591e0_0 .net "in_a", 0 0, L_0x5c7c3315b980;  alias, 1 drivers
v0x5c7c330592d0_0 .net "in_b", 0 0, L_0x5c7c3315b980;  alias, 1 drivers
v0x5c7c330593c0_0 .net "out", 0 0, L_0x5c7c3315ba30;  alias, 1 drivers
S_0x5c7c33079a60 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330583d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3307aa90_0 .net "in_a", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
v0x5c7c3307ab30_0 .net "in_b", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
v0x5c7c3307abf0_0 .net "out", 0 0, L_0x5c7c3315bd50;  alias, 1 drivers
v0x5c7c3307ad10_0 .net "temp_out", 0 0, L_0x5c7c3315bca0;  1 drivers
S_0x5c7c33079c40 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33079a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315bca0 .functor NAND 1, L_0x5c7c3315b8d0, L_0x5c7c3315b8d0, C4<1>, C4<1>;
v0x5c7c33079eb0_0 .net "in_a", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
v0x5c7c33079f70_0 .net "in_b", 0 0, L_0x5c7c3315b8d0;  alias, 1 drivers
v0x5c7c3307a0c0_0 .net "out", 0 0, L_0x5c7c3315bca0;  alias, 1 drivers
S_0x5c7c3307a1c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33079a60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3307a8e0_0 .net "in_a", 0 0, L_0x5c7c3315bca0;  alias, 1 drivers
v0x5c7c3307a980_0 .net "out", 0 0, L_0x5c7c3315bd50;  alias, 1 drivers
S_0x5c7c3307a390 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3307a1c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315bd50 .functor NAND 1, L_0x5c7c3315bca0, L_0x5c7c3315bca0, C4<1>, C4<1>;
v0x5c7c3307a600_0 .net "in_a", 0 0, L_0x5c7c3315bca0;  alias, 1 drivers
v0x5c7c3307a6f0_0 .net "in_b", 0 0, L_0x5c7c3315bca0;  alias, 1 drivers
v0x5c7c3307a7e0_0 .net "out", 0 0, L_0x5c7c3315bd50;  alias, 1 drivers
S_0x5c7c3307ae80 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330583d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3307bec0_0 .net "in_a", 0 0, L_0x5c7c3315bae0;  alias, 1 drivers
v0x5c7c3307bf90_0 .net "in_b", 0 0, L_0x5c7c3315be00;  alias, 1 drivers
v0x5c7c3307c060_0 .net "out", 0 0, L_0x5c7c3315c070;  alias, 1 drivers
v0x5c7c3307c180_0 .net "temp_out", 0 0, L_0x5c7c3315bfc0;  1 drivers
S_0x5c7c3307b060 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3307ae80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315bfc0 .functor NAND 1, L_0x5c7c3315bae0, L_0x5c7c3315be00, C4<1>, C4<1>;
v0x5c7c3307b2b0_0 .net "in_a", 0 0, L_0x5c7c3315bae0;  alias, 1 drivers
v0x5c7c3307b390_0 .net "in_b", 0 0, L_0x5c7c3315be00;  alias, 1 drivers
v0x5c7c3307b450_0 .net "out", 0 0, L_0x5c7c3315bfc0;  alias, 1 drivers
S_0x5c7c3307b5a0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3307ae80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3307bd10_0 .net "in_a", 0 0, L_0x5c7c3315bfc0;  alias, 1 drivers
v0x5c7c3307bdb0_0 .net "out", 0 0, L_0x5c7c3315c070;  alias, 1 drivers
S_0x5c7c3307b7c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3307b5a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c070 .functor NAND 1, L_0x5c7c3315bfc0, L_0x5c7c3315bfc0, C4<1>, C4<1>;
v0x5c7c3307ba30_0 .net "in_a", 0 0, L_0x5c7c3315bfc0;  alias, 1 drivers
v0x5c7c3307bb20_0 .net "in_b", 0 0, L_0x5c7c3315bfc0;  alias, 1 drivers
v0x5c7c3307bc10_0 .net "out", 0 0, L_0x5c7c3315c070;  alias, 1 drivers
S_0x5c7c3307c2d0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330583d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3307ca00_0 .net "in_a", 0 0, L_0x5c7c3315ba30;  alias, 1 drivers
v0x5c7c3307caa0_0 .net "out", 0 0, L_0x5c7c3315bae0;  alias, 1 drivers
S_0x5c7c3307c4a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3307c2d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315bae0 .functor NAND 1, L_0x5c7c3315ba30, L_0x5c7c3315ba30, C4<1>, C4<1>;
v0x5c7c3307c710_0 .net "in_a", 0 0, L_0x5c7c3315ba30;  alias, 1 drivers
v0x5c7c3307c7d0_0 .net "in_b", 0 0, L_0x5c7c3315ba30;  alias, 1 drivers
v0x5c7c3307c920_0 .net "out", 0 0, L_0x5c7c3315bae0;  alias, 1 drivers
S_0x5c7c3307cba0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330583d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3307d370_0 .net "in_a", 0 0, L_0x5c7c3315bd50;  alias, 1 drivers
v0x5c7c3307d410_0 .net "out", 0 0, L_0x5c7c3315be00;  alias, 1 drivers
S_0x5c7c3307ce10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3307cba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315be00 .functor NAND 1, L_0x5c7c3315bd50, L_0x5c7c3315bd50, C4<1>, C4<1>;
v0x5c7c3307d080_0 .net "in_a", 0 0, L_0x5c7c3315bd50;  alias, 1 drivers
v0x5c7c3307d140_0 .net "in_b", 0 0, L_0x5c7c3315bd50;  alias, 1 drivers
v0x5c7c3307d290_0 .net "out", 0 0, L_0x5c7c3315be00;  alias, 1 drivers
S_0x5c7c3307d510 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330583d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3307dcb0_0 .net "in_a", 0 0, L_0x5c7c3315c070;  alias, 1 drivers
v0x5c7c3307dd50_0 .net "out", 0 0, L_0x5c7c3315c120;  alias, 1 drivers
S_0x5c7c3307d730 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3307d510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c120 .functor NAND 1, L_0x5c7c3315c070, L_0x5c7c3315c070, C4<1>, C4<1>;
v0x5c7c3307d9a0_0 .net "in_a", 0 0, L_0x5c7c3315c070;  alias, 1 drivers
v0x5c7c3307da60_0 .net "in_b", 0 0, L_0x5c7c3315c070;  alias, 1 drivers
v0x5c7c3307dbb0_0 .net "out", 0 0, L_0x5c7c3315c120;  alias, 1 drivers
S_0x5c7c3307ecf0 .scope module, "mux_gate1" "Mux" 15 8, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330880d0_0 .net "in_a", 0 0, L_0x5c7c3315d110;  1 drivers
v0x5c7c33088170_0 .net "in_b", 0 0, L_0x5c7c3315d1b0;  1 drivers
v0x5c7c33088280_0 .net "out", 0 0, L_0x5c7c3315cf50;  1 drivers
v0x5c7c33088320_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330883c0_0 .net "sel_out", 0 0, L_0x5c7c3315c440;  1 drivers
v0x5c7c33088540_0 .net "temp_a_out", 0 0, L_0x5c7c3315c5a0;  1 drivers
v0x5c7c330886f0_0 .net "temp_b_out", 0 0, L_0x5c7c3315c700;  1 drivers
S_0x5c7c3307ef10 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c3307ecf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3307ff50_0 .net "in_a", 0 0, L_0x5c7c3315d110;  alias, 1 drivers
v0x5c7c33080020_0 .net "in_b", 0 0, L_0x5c7c3315c440;  alias, 1 drivers
v0x5c7c330800f0_0 .net "out", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
v0x5c7c33080210_0 .net "temp_out", 0 0, L_0x5c7c3315c4f0;  1 drivers
S_0x5c7c3307f160 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3307ef10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c4f0 .functor NAND 1, L_0x5c7c3315d110, L_0x5c7c3315c440, C4<1>, C4<1>;
v0x5c7c3307f3d0_0 .net "in_a", 0 0, L_0x5c7c3315d110;  alias, 1 drivers
v0x5c7c3307f4b0_0 .net "in_b", 0 0, L_0x5c7c3315c440;  alias, 1 drivers
v0x5c7c3307f570_0 .net "out", 0 0, L_0x5c7c3315c4f0;  alias, 1 drivers
S_0x5c7c3307f690 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3307ef10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3307fdd0_0 .net "in_a", 0 0, L_0x5c7c3315c4f0;  alias, 1 drivers
v0x5c7c3307fe70_0 .net "out", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
S_0x5c7c3307f8b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3307f690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c5a0 .functor NAND 1, L_0x5c7c3315c4f0, L_0x5c7c3315c4f0, C4<1>, C4<1>;
v0x5c7c3307fb20_0 .net "in_a", 0 0, L_0x5c7c3315c4f0;  alias, 1 drivers
v0x5c7c3307fbe0_0 .net "in_b", 0 0, L_0x5c7c3315c4f0;  alias, 1 drivers
v0x5c7c3307fcd0_0 .net "out", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
S_0x5c7c330802d0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c3307ecf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330812e0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33081380_0 .net "in_b", 0 0, L_0x5c7c3315d1b0;  alias, 1 drivers
v0x5c7c33081470_0 .net "out", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
v0x5c7c33081590_0 .net "temp_out", 0 0, L_0x5c7c3315c650;  1 drivers
S_0x5c7c330804b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330802d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c650 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c3315d1b0, C4<1>, C4<1>;
v0x5c7c33080720_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330807e0_0 .net "in_b", 0 0, L_0x5c7c3315d1b0;  alias, 1 drivers
v0x5c7c330808a0_0 .net "out", 0 0, L_0x5c7c3315c650;  alias, 1 drivers
S_0x5c7c330809c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330802d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33081130_0 .net "in_a", 0 0, L_0x5c7c3315c650;  alias, 1 drivers
v0x5c7c330811d0_0 .net "out", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
S_0x5c7c33080be0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330809c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c700 .functor NAND 1, L_0x5c7c3315c650, L_0x5c7c3315c650, C4<1>, C4<1>;
v0x5c7c33080e50_0 .net "in_a", 0 0, L_0x5c7c3315c650;  alias, 1 drivers
v0x5c7c33080f40_0 .net "in_b", 0 0, L_0x5c7c3315c650;  alias, 1 drivers
v0x5c7c33081030_0 .net "out", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
S_0x5c7c33081650 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c3307ecf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33081e60_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33081f00_0 .net "out", 0 0, L_0x5c7c3315c440;  alias, 1 drivers
S_0x5c7c33081820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33081650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c440 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c33081a70_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33081c40_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33081d00_0 .net "out", 0 0, L_0x5c7c3315c440;  alias, 1 drivers
S_0x5c7c33082000 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c3307ecf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33087a20_0 .net "branch1_out", 0 0, L_0x5c7c3315c910;  1 drivers
v0x5c7c33087b50_0 .net "branch2_out", 0 0, L_0x5c7c3315cc30;  1 drivers
v0x5c7c33087ca0_0 .net "in_a", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
v0x5c7c33087d70_0 .net "in_b", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
v0x5c7c33087e10_0 .net "out", 0 0, L_0x5c7c3315cf50;  alias, 1 drivers
v0x5c7c33087eb0_0 .net "temp1_out", 0 0, L_0x5c7c3315c860;  1 drivers
v0x5c7c33087f50_0 .net "temp2_out", 0 0, L_0x5c7c3315cb80;  1 drivers
v0x5c7c33087ff0_0 .net "temp3_out", 0 0, L_0x5c7c3315cea0;  1 drivers
S_0x5c7c33082230 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33082000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33083260_0 .net "in_a", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
v0x5c7c33083300_0 .net "in_b", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
v0x5c7c330833c0_0 .net "out", 0 0, L_0x5c7c3315c860;  alias, 1 drivers
v0x5c7c330834e0_0 .net "temp_out", 0 0, L_0x5c7c3315c7b0;  1 drivers
S_0x5c7c330824a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33082230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c7b0 .functor NAND 1, L_0x5c7c3315c5a0, L_0x5c7c3315c5a0, C4<1>, C4<1>;
v0x5c7c33082710_0 .net "in_a", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
v0x5c7c330827d0_0 .net "in_b", 0 0, L_0x5c7c3315c5a0;  alias, 1 drivers
v0x5c7c33082890_0 .net "out", 0 0, L_0x5c7c3315c7b0;  alias, 1 drivers
S_0x5c7c33082990 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33082230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330830b0_0 .net "in_a", 0 0, L_0x5c7c3315c7b0;  alias, 1 drivers
v0x5c7c33083150_0 .net "out", 0 0, L_0x5c7c3315c860;  alias, 1 drivers
S_0x5c7c33082b60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33082990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c860 .functor NAND 1, L_0x5c7c3315c7b0, L_0x5c7c3315c7b0, C4<1>, C4<1>;
v0x5c7c33082dd0_0 .net "in_a", 0 0, L_0x5c7c3315c7b0;  alias, 1 drivers
v0x5c7c33082ec0_0 .net "in_b", 0 0, L_0x5c7c3315c7b0;  alias, 1 drivers
v0x5c7c33082fb0_0 .net "out", 0 0, L_0x5c7c3315c860;  alias, 1 drivers
S_0x5c7c33083650 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33082000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33084680_0 .net "in_a", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
v0x5c7c33084720_0 .net "in_b", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
v0x5c7c330847e0_0 .net "out", 0 0, L_0x5c7c3315cb80;  alias, 1 drivers
v0x5c7c33084900_0 .net "temp_out", 0 0, L_0x5c7c3315cad0;  1 drivers
S_0x5c7c33083830 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33083650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315cad0 .functor NAND 1, L_0x5c7c3315c700, L_0x5c7c3315c700, C4<1>, C4<1>;
v0x5c7c33083aa0_0 .net "in_a", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
v0x5c7c33083b60_0 .net "in_b", 0 0, L_0x5c7c3315c700;  alias, 1 drivers
v0x5c7c33083cb0_0 .net "out", 0 0, L_0x5c7c3315cad0;  alias, 1 drivers
S_0x5c7c33083db0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33083650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330844d0_0 .net "in_a", 0 0, L_0x5c7c3315cad0;  alias, 1 drivers
v0x5c7c33084570_0 .net "out", 0 0, L_0x5c7c3315cb80;  alias, 1 drivers
S_0x5c7c33083f80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33083db0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315cb80 .functor NAND 1, L_0x5c7c3315cad0, L_0x5c7c3315cad0, C4<1>, C4<1>;
v0x5c7c330841f0_0 .net "in_a", 0 0, L_0x5c7c3315cad0;  alias, 1 drivers
v0x5c7c330842e0_0 .net "in_b", 0 0, L_0x5c7c3315cad0;  alias, 1 drivers
v0x5c7c330843d0_0 .net "out", 0 0, L_0x5c7c3315cb80;  alias, 1 drivers
S_0x5c7c33084a70 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33082000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33085ab0_0 .net "in_a", 0 0, L_0x5c7c3315c910;  alias, 1 drivers
v0x5c7c33085b80_0 .net "in_b", 0 0, L_0x5c7c3315cc30;  alias, 1 drivers
v0x5c7c33085c50_0 .net "out", 0 0, L_0x5c7c3315cea0;  alias, 1 drivers
v0x5c7c33085d70_0 .net "temp_out", 0 0, L_0x5c7c3315cdf0;  1 drivers
S_0x5c7c33084c50 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33084a70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315cdf0 .functor NAND 1, L_0x5c7c3315c910, L_0x5c7c3315cc30, C4<1>, C4<1>;
v0x5c7c33084ea0_0 .net "in_a", 0 0, L_0x5c7c3315c910;  alias, 1 drivers
v0x5c7c33084f80_0 .net "in_b", 0 0, L_0x5c7c3315cc30;  alias, 1 drivers
v0x5c7c33085040_0 .net "out", 0 0, L_0x5c7c3315cdf0;  alias, 1 drivers
S_0x5c7c33085190 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33084a70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33085900_0 .net "in_a", 0 0, L_0x5c7c3315cdf0;  alias, 1 drivers
v0x5c7c330859a0_0 .net "out", 0 0, L_0x5c7c3315cea0;  alias, 1 drivers
S_0x5c7c330853b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33085190;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315cea0 .functor NAND 1, L_0x5c7c3315cdf0, L_0x5c7c3315cdf0, C4<1>, C4<1>;
v0x5c7c33085620_0 .net "in_a", 0 0, L_0x5c7c3315cdf0;  alias, 1 drivers
v0x5c7c33085710_0 .net "in_b", 0 0, L_0x5c7c3315cdf0;  alias, 1 drivers
v0x5c7c33085800_0 .net "out", 0 0, L_0x5c7c3315cea0;  alias, 1 drivers
S_0x5c7c33085ec0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33082000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330865f0_0 .net "in_a", 0 0, L_0x5c7c3315c860;  alias, 1 drivers
v0x5c7c33086690_0 .net "out", 0 0, L_0x5c7c3315c910;  alias, 1 drivers
S_0x5c7c33086090 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33085ec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315c910 .functor NAND 1, L_0x5c7c3315c860, L_0x5c7c3315c860, C4<1>, C4<1>;
v0x5c7c33086300_0 .net "in_a", 0 0, L_0x5c7c3315c860;  alias, 1 drivers
v0x5c7c330863c0_0 .net "in_b", 0 0, L_0x5c7c3315c860;  alias, 1 drivers
v0x5c7c33086510_0 .net "out", 0 0, L_0x5c7c3315c910;  alias, 1 drivers
S_0x5c7c33086790 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33082000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33086f60_0 .net "in_a", 0 0, L_0x5c7c3315cb80;  alias, 1 drivers
v0x5c7c33087000_0 .net "out", 0 0, L_0x5c7c3315cc30;  alias, 1 drivers
S_0x5c7c33086a00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33086790;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315cc30 .functor NAND 1, L_0x5c7c3315cb80, L_0x5c7c3315cb80, C4<1>, C4<1>;
v0x5c7c33086c70_0 .net "in_a", 0 0, L_0x5c7c3315cb80;  alias, 1 drivers
v0x5c7c33086d30_0 .net "in_b", 0 0, L_0x5c7c3315cb80;  alias, 1 drivers
v0x5c7c33086e80_0 .net "out", 0 0, L_0x5c7c3315cc30;  alias, 1 drivers
S_0x5c7c33087100 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33082000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330878a0_0 .net "in_a", 0 0, L_0x5c7c3315cea0;  alias, 1 drivers
v0x5c7c33087940_0 .net "out", 0 0, L_0x5c7c3315cf50;  alias, 1 drivers
S_0x5c7c33087320 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33087100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315cf50 .functor NAND 1, L_0x5c7c3315cea0, L_0x5c7c3315cea0, C4<1>, C4<1>;
v0x5c7c33087590_0 .net "in_a", 0 0, L_0x5c7c3315cea0;  alias, 1 drivers
v0x5c7c33087650_0 .net "in_b", 0 0, L_0x5c7c3315cea0;  alias, 1 drivers
v0x5c7c330877a0_0 .net "out", 0 0, L_0x5c7c3315cf50;  alias, 1 drivers
S_0x5c7c330888e0 .scope module, "mux_gate10" "Mux" 15 17, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33091c50_0 .net "in_a", 0 0, L_0x5c7c33163870;  1 drivers
v0x5c7c33091cf0_0 .net "in_b", 0 0, L_0x5c7c33165be0;  1 drivers
v0x5c7c33091e00_0 .net "out", 0 0, L_0x5c7c33165a60;  1 drivers
v0x5c7c33091ea0_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33091f40_0 .net "sel_out", 0 0, L_0x5c7c331647d0;  1 drivers
v0x5c7c330920c0_0 .net "temp_a_out", 0 0, L_0x5c7c330d9570;  1 drivers
v0x5c7c33092160_0 .net "temp_b_out", 0 0, L_0x5c7c330d96d0;  1 drivers
S_0x5c7c33088ae0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330888e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33089b50_0 .net "in_a", 0 0, L_0x5c7c33163870;  alias, 1 drivers
v0x5c7c33089c20_0 .net "in_b", 0 0, L_0x5c7c331647d0;  alias, 1 drivers
v0x5c7c33089cf0_0 .net "out", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
v0x5c7c33089e10_0 .net "temp_out", 0 0, L_0x5c7c330d94c0;  1 drivers
S_0x5c7c33088d30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33088ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d94c0 .functor NAND 1, L_0x5c7c33163870, L_0x5c7c331647d0, C4<1>, C4<1>;
v0x5c7c33088fa0_0 .net "in_a", 0 0, L_0x5c7c33163870;  alias, 1 drivers
v0x5c7c33089080_0 .net "in_b", 0 0, L_0x5c7c331647d0;  alias, 1 drivers
v0x5c7c33089140_0 .net "out", 0 0, L_0x5c7c330d94c0;  alias, 1 drivers
S_0x5c7c33089260 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33088ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330899a0_0 .net "in_a", 0 0, L_0x5c7c330d94c0;  alias, 1 drivers
v0x5c7c33089a40_0 .net "out", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
S_0x5c7c33089480 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33089260;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9570 .functor NAND 1, L_0x5c7c330d94c0, L_0x5c7c330d94c0, C4<1>, C4<1>;
v0x5c7c330896f0_0 .net "in_a", 0 0, L_0x5c7c330d94c0;  alias, 1 drivers
v0x5c7c330897b0_0 .net "in_b", 0 0, L_0x5c7c330d94c0;  alias, 1 drivers
v0x5c7c330898a0_0 .net "out", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
S_0x5c7c33089ed0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330888e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3308aee0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3308af80_0 .net "in_b", 0 0, L_0x5c7c33165be0;  alias, 1 drivers
v0x5c7c3308b070_0 .net "out", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
v0x5c7c3308b190_0 .net "temp_out", 0 0, L_0x5c7c330d9620;  1 drivers
S_0x5c7c3308a0b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33089ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9620 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33165be0, C4<1>, C4<1>;
v0x5c7c3308a320_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3308a3e0_0 .net "in_b", 0 0, L_0x5c7c33165be0;  alias, 1 drivers
v0x5c7c3308a4a0_0 .net "out", 0 0, L_0x5c7c330d9620;  alias, 1 drivers
S_0x5c7c3308a5c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33089ed0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3308ad30_0 .net "in_a", 0 0, L_0x5c7c330d9620;  alias, 1 drivers
v0x5c7c3308add0_0 .net "out", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
S_0x5c7c3308a7e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3308a5c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d96d0 .functor NAND 1, L_0x5c7c330d9620, L_0x5c7c330d9620, C4<1>, C4<1>;
v0x5c7c3308aa50_0 .net "in_a", 0 0, L_0x5c7c330d9620;  alias, 1 drivers
v0x5c7c3308ab40_0 .net "in_b", 0 0, L_0x5c7c330d9620;  alias, 1 drivers
v0x5c7c3308ac30_0 .net "out", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
S_0x5c7c3308b250 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330888e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3308b950_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3308b9f0_0 .net "out", 0 0, L_0x5c7c331647d0;  alias, 1 drivers
S_0x5c7c3308b420 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3308b250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331647d0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c3308b670_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3308b730_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3308b7f0_0 .net "out", 0 0, L_0x5c7c331647d0;  alias, 1 drivers
S_0x5c7c3308baf0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330888e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330915a0_0 .net "branch1_out", 0 0, L_0x5c7c330d98e0;  1 drivers
v0x5c7c330916d0_0 .net "branch2_out", 0 0, L_0x5c7c330d9c00;  1 drivers
v0x5c7c33091820_0 .net "in_a", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
v0x5c7c330918f0_0 .net "in_b", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
v0x5c7c33091990_0 .net "out", 0 0, L_0x5c7c33165a60;  alias, 1 drivers
v0x5c7c33091a30_0 .net "temp1_out", 0 0, L_0x5c7c330d9830;  1 drivers
v0x5c7c33091ad0_0 .net "temp2_out", 0 0, L_0x5c7c330d9b50;  1 drivers
v0x5c7c33091b70_0 .net "temp3_out", 0 0, L_0x5c7c331659f0;  1 drivers
S_0x5c7c3308bd20 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c3308baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3308cde0_0 .net "in_a", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
v0x5c7c3308ce80_0 .net "in_b", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
v0x5c7c3308cf40_0 .net "out", 0 0, L_0x5c7c330d9830;  alias, 1 drivers
v0x5c7c3308d060_0 .net "temp_out", 0 0, L_0x5c7c330d9780;  1 drivers
S_0x5c7c3308bf90 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3308bd20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9780 .functor NAND 1, L_0x5c7c330d9570, L_0x5c7c330d9570, C4<1>, C4<1>;
v0x5c7c3308c200_0 .net "in_a", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
v0x5c7c3308c2c0_0 .net "in_b", 0 0, L_0x5c7c330d9570;  alias, 1 drivers
v0x5c7c3308c410_0 .net "out", 0 0, L_0x5c7c330d9780;  alias, 1 drivers
S_0x5c7c3308c510 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3308bd20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3308cc30_0 .net "in_a", 0 0, L_0x5c7c330d9780;  alias, 1 drivers
v0x5c7c3308ccd0_0 .net "out", 0 0, L_0x5c7c330d9830;  alias, 1 drivers
S_0x5c7c3308c6e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3308c510;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9830 .functor NAND 1, L_0x5c7c330d9780, L_0x5c7c330d9780, C4<1>, C4<1>;
v0x5c7c3308c950_0 .net "in_a", 0 0, L_0x5c7c330d9780;  alias, 1 drivers
v0x5c7c3308ca40_0 .net "in_b", 0 0, L_0x5c7c330d9780;  alias, 1 drivers
v0x5c7c3308cb30_0 .net "out", 0 0, L_0x5c7c330d9830;  alias, 1 drivers
S_0x5c7c3308d1d0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c3308baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3308e200_0 .net "in_a", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
v0x5c7c3308e2a0_0 .net "in_b", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
v0x5c7c3308e360_0 .net "out", 0 0, L_0x5c7c330d9b50;  alias, 1 drivers
v0x5c7c3308e480_0 .net "temp_out", 0 0, L_0x5c7c330d9aa0;  1 drivers
S_0x5c7c3308d3b0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3308d1d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9aa0 .functor NAND 1, L_0x5c7c330d96d0, L_0x5c7c330d96d0, C4<1>, C4<1>;
v0x5c7c3308d620_0 .net "in_a", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
v0x5c7c3308d6e0_0 .net "in_b", 0 0, L_0x5c7c330d96d0;  alias, 1 drivers
v0x5c7c3308d830_0 .net "out", 0 0, L_0x5c7c330d9aa0;  alias, 1 drivers
S_0x5c7c3308d930 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3308d1d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3308e050_0 .net "in_a", 0 0, L_0x5c7c330d9aa0;  alias, 1 drivers
v0x5c7c3308e0f0_0 .net "out", 0 0, L_0x5c7c330d9b50;  alias, 1 drivers
S_0x5c7c3308db00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3308d930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9b50 .functor NAND 1, L_0x5c7c330d9aa0, L_0x5c7c330d9aa0, C4<1>, C4<1>;
v0x5c7c3308dd70_0 .net "in_a", 0 0, L_0x5c7c330d9aa0;  alias, 1 drivers
v0x5c7c3308de60_0 .net "in_b", 0 0, L_0x5c7c330d9aa0;  alias, 1 drivers
v0x5c7c3308df50_0 .net "out", 0 0, L_0x5c7c330d9b50;  alias, 1 drivers
S_0x5c7c3308e5f0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c3308baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3308f630_0 .net "in_a", 0 0, L_0x5c7c330d98e0;  alias, 1 drivers
v0x5c7c3308f700_0 .net "in_b", 0 0, L_0x5c7c330d9c00;  alias, 1 drivers
v0x5c7c3308f7d0_0 .net "out", 0 0, L_0x5c7c331659f0;  alias, 1 drivers
v0x5c7c3308f8f0_0 .net "temp_out", 0 0, L_0x5c7c33165980;  1 drivers
S_0x5c7c3308e7d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3308e5f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165980 .functor NAND 1, L_0x5c7c330d98e0, L_0x5c7c330d9c00, C4<1>, C4<1>;
v0x5c7c3308ea20_0 .net "in_a", 0 0, L_0x5c7c330d98e0;  alias, 1 drivers
v0x5c7c3308eb00_0 .net "in_b", 0 0, L_0x5c7c330d9c00;  alias, 1 drivers
v0x5c7c3308ebc0_0 .net "out", 0 0, L_0x5c7c33165980;  alias, 1 drivers
S_0x5c7c3308ed10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3308e5f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3308f480_0 .net "in_a", 0 0, L_0x5c7c33165980;  alias, 1 drivers
v0x5c7c3308f520_0 .net "out", 0 0, L_0x5c7c331659f0;  alias, 1 drivers
S_0x5c7c3308ef30 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3308ed10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331659f0 .functor NAND 1, L_0x5c7c33165980, L_0x5c7c33165980, C4<1>, C4<1>;
v0x5c7c3308f1a0_0 .net "in_a", 0 0, L_0x5c7c33165980;  alias, 1 drivers
v0x5c7c3308f290_0 .net "in_b", 0 0, L_0x5c7c33165980;  alias, 1 drivers
v0x5c7c3308f380_0 .net "out", 0 0, L_0x5c7c331659f0;  alias, 1 drivers
S_0x5c7c3308fa40 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c3308baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33090170_0 .net "in_a", 0 0, L_0x5c7c330d9830;  alias, 1 drivers
v0x5c7c33090210_0 .net "out", 0 0, L_0x5c7c330d98e0;  alias, 1 drivers
S_0x5c7c3308fc10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3308fa40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d98e0 .functor NAND 1, L_0x5c7c330d9830, L_0x5c7c330d9830, C4<1>, C4<1>;
v0x5c7c3308fe80_0 .net "in_a", 0 0, L_0x5c7c330d9830;  alias, 1 drivers
v0x5c7c3308ff40_0 .net "in_b", 0 0, L_0x5c7c330d9830;  alias, 1 drivers
v0x5c7c33090090_0 .net "out", 0 0, L_0x5c7c330d98e0;  alias, 1 drivers
S_0x5c7c33090310 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c3308baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33090ae0_0 .net "in_a", 0 0, L_0x5c7c330d9b50;  alias, 1 drivers
v0x5c7c33090b80_0 .net "out", 0 0, L_0x5c7c330d9c00;  alias, 1 drivers
S_0x5c7c33090580 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33090310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c330d9c00 .functor NAND 1, L_0x5c7c330d9b50, L_0x5c7c330d9b50, C4<1>, C4<1>;
v0x5c7c330907f0_0 .net "in_a", 0 0, L_0x5c7c330d9b50;  alias, 1 drivers
v0x5c7c330908b0_0 .net "in_b", 0 0, L_0x5c7c330d9b50;  alias, 1 drivers
v0x5c7c33090a00_0 .net "out", 0 0, L_0x5c7c330d9c00;  alias, 1 drivers
S_0x5c7c33090c80 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c3308baf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33091420_0 .net "in_a", 0 0, L_0x5c7c331659f0;  alias, 1 drivers
v0x5c7c330914c0_0 .net "out", 0 0, L_0x5c7c33165a60;  alias, 1 drivers
S_0x5c7c33090ea0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33090c80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165a60 .functor NAND 1, L_0x5c7c331659f0, L_0x5c7c331659f0, C4<1>, C4<1>;
v0x5c7c33091110_0 .net "in_a", 0 0, L_0x5c7c331659f0;  alias, 1 drivers
v0x5c7c330911d0_0 .net "in_b", 0 0, L_0x5c7c331659f0;  alias, 1 drivers
v0x5c7c33091320_0 .net "out", 0 0, L_0x5c7c33165a60;  alias, 1 drivers
S_0x5c7c33092350 .scope module, "mux_gate11" "Mux" 15 18, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c3309b6b0_0 .net "in_a", 0 0, L_0x5c7c33166690;  1 drivers
v0x5c7c3309b750_0 .net "in_b", 0 0, L_0x5c7c33166730;  1 drivers
v0x5c7c3309b860_0 .net "out", 0 0, L_0x5c7c33166510;  1 drivers
v0x5c7c3309b900_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3309b9a0_0 .net "sel_out", 0 0, L_0x5c7c33165d40;  1 drivers
v0x5c7c3309bb20_0 .net "temp_a_out", 0 0, L_0x5c7c33165e20;  1 drivers
v0x5c7c3309bcd0_0 .net "temp_b_out", 0 0, L_0x5c7c33165f00;  1 drivers
S_0x5c7c33092550 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33092350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330935b0_0 .net "in_a", 0 0, L_0x5c7c33166690;  alias, 1 drivers
v0x5c7c33093680_0 .net "in_b", 0 0, L_0x5c7c33165d40;  alias, 1 drivers
v0x5c7c33093750_0 .net "out", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
v0x5c7c33093870_0 .net "temp_out", 0 0, L_0x5c7c33165db0;  1 drivers
S_0x5c7c330927c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33092550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165db0 .functor NAND 1, L_0x5c7c33166690, L_0x5c7c33165d40, C4<1>, C4<1>;
v0x5c7c33092a30_0 .net "in_a", 0 0, L_0x5c7c33166690;  alias, 1 drivers
v0x5c7c33092b10_0 .net "in_b", 0 0, L_0x5c7c33165d40;  alias, 1 drivers
v0x5c7c33092bd0_0 .net "out", 0 0, L_0x5c7c33165db0;  alias, 1 drivers
S_0x5c7c33092cf0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33092550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33093430_0 .net "in_a", 0 0, L_0x5c7c33165db0;  alias, 1 drivers
v0x5c7c330934d0_0 .net "out", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
S_0x5c7c33092f10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33092cf0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165e20 .functor NAND 1, L_0x5c7c33165db0, L_0x5c7c33165db0, C4<1>, C4<1>;
v0x5c7c33093180_0 .net "in_a", 0 0, L_0x5c7c33165db0;  alias, 1 drivers
v0x5c7c33093240_0 .net "in_b", 0 0, L_0x5c7c33165db0;  alias, 1 drivers
v0x5c7c33093330_0 .net "out", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
S_0x5c7c33093930 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33092350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33094940_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330949e0_0 .net "in_b", 0 0, L_0x5c7c33166730;  alias, 1 drivers
v0x5c7c33094ad0_0 .net "out", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
v0x5c7c33094bf0_0 .net "temp_out", 0 0, L_0x5c7c33165e90;  1 drivers
S_0x5c7c33093b10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33093930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165e90 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33166730, C4<1>, C4<1>;
v0x5c7c33093d80_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33093e40_0 .net "in_b", 0 0, L_0x5c7c33166730;  alias, 1 drivers
v0x5c7c33093f00_0 .net "out", 0 0, L_0x5c7c33165e90;  alias, 1 drivers
S_0x5c7c33094020 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33093930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33094790_0 .net "in_a", 0 0, L_0x5c7c33165e90;  alias, 1 drivers
v0x5c7c33094830_0 .net "out", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
S_0x5c7c33094240 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33094020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165f00 .functor NAND 1, L_0x5c7c33165e90, L_0x5c7c33165e90, C4<1>, C4<1>;
v0x5c7c330944b0_0 .net "in_a", 0 0, L_0x5c7c33165e90;  alias, 1 drivers
v0x5c7c330945a0_0 .net "in_b", 0 0, L_0x5c7c33165e90;  alias, 1 drivers
v0x5c7c33094690_0 .net "out", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
S_0x5c7c33094cb0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33092350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330953b0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33095450_0 .net "out", 0 0, L_0x5c7c33165d40;  alias, 1 drivers
S_0x5c7c33094e80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33094cb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165d40 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330950d0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33095190_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33095250_0 .net "out", 0 0, L_0x5c7c33165d40;  alias, 1 drivers
S_0x5c7c33095550 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33092350;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3309b000_0 .net "branch1_out", 0 0, L_0x5c7c33166050;  1 drivers
v0x5c7c3309b130_0 .net "branch2_out", 0 0, L_0x5c7c331662b0;  1 drivers
v0x5c7c3309b280_0 .net "in_a", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
v0x5c7c3309b350_0 .net "in_b", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
v0x5c7c3309b3f0_0 .net "out", 0 0, L_0x5c7c33166510;  alias, 1 drivers
v0x5c7c3309b490_0 .net "temp1_out", 0 0, L_0x5c7c33165fe0;  1 drivers
v0x5c7c3309b530_0 .net "temp2_out", 0 0, L_0x5c7c33166240;  1 drivers
v0x5c7c3309b5d0_0 .net "temp3_out", 0 0, L_0x5c7c331664a0;  1 drivers
S_0x5c7c33095780 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33095550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33096840_0 .net "in_a", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
v0x5c7c330968e0_0 .net "in_b", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
v0x5c7c330969a0_0 .net "out", 0 0, L_0x5c7c33165fe0;  alias, 1 drivers
v0x5c7c33096ac0_0 .net "temp_out", 0 0, L_0x5c7c33165f70;  1 drivers
S_0x5c7c330959f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33095780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165f70 .functor NAND 1, L_0x5c7c33165e20, L_0x5c7c33165e20, C4<1>, C4<1>;
v0x5c7c33095c60_0 .net "in_a", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
v0x5c7c33095d20_0 .net "in_b", 0 0, L_0x5c7c33165e20;  alias, 1 drivers
v0x5c7c33095e70_0 .net "out", 0 0, L_0x5c7c33165f70;  alias, 1 drivers
S_0x5c7c33095f70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33095780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33096690_0 .net "in_a", 0 0, L_0x5c7c33165f70;  alias, 1 drivers
v0x5c7c33096730_0 .net "out", 0 0, L_0x5c7c33165fe0;  alias, 1 drivers
S_0x5c7c33096140 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33095f70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33165fe0 .functor NAND 1, L_0x5c7c33165f70, L_0x5c7c33165f70, C4<1>, C4<1>;
v0x5c7c330963b0_0 .net "in_a", 0 0, L_0x5c7c33165f70;  alias, 1 drivers
v0x5c7c330964a0_0 .net "in_b", 0 0, L_0x5c7c33165f70;  alias, 1 drivers
v0x5c7c33096590_0 .net "out", 0 0, L_0x5c7c33165fe0;  alias, 1 drivers
S_0x5c7c33096c30 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33095550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33097c60_0 .net "in_a", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
v0x5c7c33097d00_0 .net "in_b", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
v0x5c7c33097dc0_0 .net "out", 0 0, L_0x5c7c33166240;  alias, 1 drivers
v0x5c7c33097ee0_0 .net "temp_out", 0 0, L_0x5c7c331661d0;  1 drivers
S_0x5c7c33096e10 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33096c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331661d0 .functor NAND 1, L_0x5c7c33165f00, L_0x5c7c33165f00, C4<1>, C4<1>;
v0x5c7c33097080_0 .net "in_a", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
v0x5c7c33097140_0 .net "in_b", 0 0, L_0x5c7c33165f00;  alias, 1 drivers
v0x5c7c33097290_0 .net "out", 0 0, L_0x5c7c331661d0;  alias, 1 drivers
S_0x5c7c33097390 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33096c30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33097ab0_0 .net "in_a", 0 0, L_0x5c7c331661d0;  alias, 1 drivers
v0x5c7c33097b50_0 .net "out", 0 0, L_0x5c7c33166240;  alias, 1 drivers
S_0x5c7c33097560 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33097390;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166240 .functor NAND 1, L_0x5c7c331661d0, L_0x5c7c331661d0, C4<1>, C4<1>;
v0x5c7c330977d0_0 .net "in_a", 0 0, L_0x5c7c331661d0;  alias, 1 drivers
v0x5c7c330978c0_0 .net "in_b", 0 0, L_0x5c7c331661d0;  alias, 1 drivers
v0x5c7c330979b0_0 .net "out", 0 0, L_0x5c7c33166240;  alias, 1 drivers
S_0x5c7c33098050 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33095550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33099090_0 .net "in_a", 0 0, L_0x5c7c33166050;  alias, 1 drivers
v0x5c7c33099160_0 .net "in_b", 0 0, L_0x5c7c331662b0;  alias, 1 drivers
v0x5c7c33099230_0 .net "out", 0 0, L_0x5c7c331664a0;  alias, 1 drivers
v0x5c7c33099350_0 .net "temp_out", 0 0, L_0x5c7c33166430;  1 drivers
S_0x5c7c33098230 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33098050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166430 .functor NAND 1, L_0x5c7c33166050, L_0x5c7c331662b0, C4<1>, C4<1>;
v0x5c7c33098480_0 .net "in_a", 0 0, L_0x5c7c33166050;  alias, 1 drivers
v0x5c7c33098560_0 .net "in_b", 0 0, L_0x5c7c331662b0;  alias, 1 drivers
v0x5c7c33098620_0 .net "out", 0 0, L_0x5c7c33166430;  alias, 1 drivers
S_0x5c7c33098770 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33098050;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33098ee0_0 .net "in_a", 0 0, L_0x5c7c33166430;  alias, 1 drivers
v0x5c7c33098f80_0 .net "out", 0 0, L_0x5c7c331664a0;  alias, 1 drivers
S_0x5c7c33098990 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33098770;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331664a0 .functor NAND 1, L_0x5c7c33166430, L_0x5c7c33166430, C4<1>, C4<1>;
v0x5c7c33098c00_0 .net "in_a", 0 0, L_0x5c7c33166430;  alias, 1 drivers
v0x5c7c33098cf0_0 .net "in_b", 0 0, L_0x5c7c33166430;  alias, 1 drivers
v0x5c7c33098de0_0 .net "out", 0 0, L_0x5c7c331664a0;  alias, 1 drivers
S_0x5c7c330994a0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33095550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33099bd0_0 .net "in_a", 0 0, L_0x5c7c33165fe0;  alias, 1 drivers
v0x5c7c33099c70_0 .net "out", 0 0, L_0x5c7c33166050;  alias, 1 drivers
S_0x5c7c33099670 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330994a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166050 .functor NAND 1, L_0x5c7c33165fe0, L_0x5c7c33165fe0, C4<1>, C4<1>;
v0x5c7c330998e0_0 .net "in_a", 0 0, L_0x5c7c33165fe0;  alias, 1 drivers
v0x5c7c330999a0_0 .net "in_b", 0 0, L_0x5c7c33165fe0;  alias, 1 drivers
v0x5c7c33099af0_0 .net "out", 0 0, L_0x5c7c33166050;  alias, 1 drivers
S_0x5c7c33099d70 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33095550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3309a540_0 .net "in_a", 0 0, L_0x5c7c33166240;  alias, 1 drivers
v0x5c7c3309a5e0_0 .net "out", 0 0, L_0x5c7c331662b0;  alias, 1 drivers
S_0x5c7c33099fe0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33099d70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331662b0 .functor NAND 1, L_0x5c7c33166240, L_0x5c7c33166240, C4<1>, C4<1>;
v0x5c7c3309a250_0 .net "in_a", 0 0, L_0x5c7c33166240;  alias, 1 drivers
v0x5c7c3309a310_0 .net "in_b", 0 0, L_0x5c7c33166240;  alias, 1 drivers
v0x5c7c3309a460_0 .net "out", 0 0, L_0x5c7c331662b0;  alias, 1 drivers
S_0x5c7c3309a6e0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33095550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3309ae80_0 .net "in_a", 0 0, L_0x5c7c331664a0;  alias, 1 drivers
v0x5c7c3309af20_0 .net "out", 0 0, L_0x5c7c33166510;  alias, 1 drivers
S_0x5c7c3309a900 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3309a6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166510 .functor NAND 1, L_0x5c7c331664a0, L_0x5c7c331664a0, C4<1>, C4<1>;
v0x5c7c3309ab70_0 .net "in_a", 0 0, L_0x5c7c331664a0;  alias, 1 drivers
v0x5c7c3309ac30_0 .net "in_b", 0 0, L_0x5c7c331664a0;  alias, 1 drivers
v0x5c7c3309ad80_0 .net "out", 0 0, L_0x5c7c33166510;  alias, 1 drivers
S_0x5c7c3309bec0 .scope module, "mux_gate12" "Mux" 15 19, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330a5240_0 .net "in_a", 0 0, L_0x5c7c331671f0;  1 drivers
v0x5c7c330a52e0_0 .net "in_b", 0 0, L_0x5c7c331674a0;  1 drivers
v0x5c7c330a53f0_0 .net "out", 0 0, L_0x5c7c33167070;  1 drivers
v0x5c7c330a5490_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330a5530_0 .net "sel_out", 0 0, L_0x5c7c331668a0;  1 drivers
v0x5c7c330a56b0_0 .net "temp_a_out", 0 0, L_0x5c7c33166980;  1 drivers
v0x5c7c330a5860_0 .net "temp_b_out", 0 0, L_0x5c7c33166a60;  1 drivers
S_0x5c7c3309c110 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c3309bec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3309d170_0 .net "in_a", 0 0, L_0x5c7c331671f0;  alias, 1 drivers
v0x5c7c3309d210_0 .net "in_b", 0 0, L_0x5c7c331668a0;  alias, 1 drivers
v0x5c7c3309d2e0_0 .net "out", 0 0, L_0x5c7c33166980;  alias, 1 drivers
v0x5c7c3309d400_0 .net "temp_out", 0 0, L_0x5c7c33166910;  1 drivers
S_0x5c7c3309c380 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3309c110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166910 .functor NAND 1, L_0x5c7c331671f0, L_0x5c7c331668a0, C4<1>, C4<1>;
v0x5c7c3309c5f0_0 .net "in_a", 0 0, L_0x5c7c331671f0;  alias, 1 drivers
v0x5c7c3309c6d0_0 .net "in_b", 0 0, L_0x5c7c331668a0;  alias, 1 drivers
v0x5c7c3309c790_0 .net "out", 0 0, L_0x5c7c33166910;  alias, 1 drivers
S_0x5c7c3309c8b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3309c110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3309cff0_0 .net "in_a", 0 0, L_0x5c7c33166910;  alias, 1 drivers
v0x5c7c3309d090_0 .net "out", 0 0, L_0x5c7c33166980;  alias, 1 drivers
S_0x5c7c3309cad0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3309c8b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166980 .functor NAND 1, L_0x5c7c33166910, L_0x5c7c33166910, C4<1>, C4<1>;
v0x5c7c3309cd40_0 .net "in_a", 0 0, L_0x5c7c33166910;  alias, 1 drivers
v0x5c7c3309ce00_0 .net "in_b", 0 0, L_0x5c7c33166910;  alias, 1 drivers
v0x5c7c3309cef0_0 .net "out", 0 0, L_0x5c7c33166980;  alias, 1 drivers
S_0x5c7c3309d4c0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c3309bec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3309e4d0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3309e570_0 .net "in_b", 0 0, L_0x5c7c331674a0;  alias, 1 drivers
v0x5c7c3309e660_0 .net "out", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
v0x5c7c3309e780_0 .net "temp_out", 0 0, L_0x5c7c331669f0;  1 drivers
S_0x5c7c3309d6a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3309d4c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331669f0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c331674a0, C4<1>, C4<1>;
v0x5c7c3309d910_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3309d9d0_0 .net "in_b", 0 0, L_0x5c7c331674a0;  alias, 1 drivers
v0x5c7c3309da90_0 .net "out", 0 0, L_0x5c7c331669f0;  alias, 1 drivers
S_0x5c7c3309dbb0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3309d4c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3309e320_0 .net "in_a", 0 0, L_0x5c7c331669f0;  alias, 1 drivers
v0x5c7c3309e3c0_0 .net "out", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
S_0x5c7c3309ddd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3309dbb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166a60 .functor NAND 1, L_0x5c7c331669f0, L_0x5c7c331669f0, C4<1>, C4<1>;
v0x5c7c3309e040_0 .net "in_a", 0 0, L_0x5c7c331669f0;  alias, 1 drivers
v0x5c7c3309e130_0 .net "in_b", 0 0, L_0x5c7c331669f0;  alias, 1 drivers
v0x5c7c3309e220_0 .net "out", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
S_0x5c7c3309e840 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c3309bec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3309ef40_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3309efe0_0 .net "out", 0 0, L_0x5c7c331668a0;  alias, 1 drivers
S_0x5c7c3309ea10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3309e840;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331668a0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c3309ec60_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3309ed20_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3309ede0_0 .net "out", 0 0, L_0x5c7c331668a0;  alias, 1 drivers
S_0x5c7c3309f0e0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c3309bec0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a4b90_0 .net "branch1_out", 0 0, L_0x5c7c33166bb0;  1 drivers
v0x5c7c330a4cc0_0 .net "branch2_out", 0 0, L_0x5c7c33166e10;  1 drivers
v0x5c7c330a4e10_0 .net "in_a", 0 0, L_0x5c7c33166980;  alias, 1 drivers
v0x5c7c330a4ee0_0 .net "in_b", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
v0x5c7c330a4f80_0 .net "out", 0 0, L_0x5c7c33167070;  alias, 1 drivers
v0x5c7c330a5020_0 .net "temp1_out", 0 0, L_0x5c7c33166b40;  1 drivers
v0x5c7c330a50c0_0 .net "temp2_out", 0 0, L_0x5c7c33166da0;  1 drivers
v0x5c7c330a5160_0 .net "temp3_out", 0 0, L_0x5c7c33167000;  1 drivers
S_0x5c7c3309f310 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c3309f0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a03d0_0 .net "in_a", 0 0, L_0x5c7c33166980;  alias, 1 drivers
v0x5c7c330a0470_0 .net "in_b", 0 0, L_0x5c7c33166980;  alias, 1 drivers
v0x5c7c330a0530_0 .net "out", 0 0, L_0x5c7c33166b40;  alias, 1 drivers
v0x5c7c330a0650_0 .net "temp_out", 0 0, L_0x5c7c33166ad0;  1 drivers
S_0x5c7c3309f580 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3309f310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166ad0 .functor NAND 1, L_0x5c7c33166980, L_0x5c7c33166980, C4<1>, C4<1>;
v0x5c7c3309f7f0_0 .net "in_a", 0 0, L_0x5c7c33166980;  alias, 1 drivers
v0x5c7c3309f8b0_0 .net "in_b", 0 0, L_0x5c7c33166980;  alias, 1 drivers
v0x5c7c3309fa00_0 .net "out", 0 0, L_0x5c7c33166ad0;  alias, 1 drivers
S_0x5c7c3309fb00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3309f310;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a0220_0 .net "in_a", 0 0, L_0x5c7c33166ad0;  alias, 1 drivers
v0x5c7c330a02c0_0 .net "out", 0 0, L_0x5c7c33166b40;  alias, 1 drivers
S_0x5c7c3309fcd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3309fb00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166b40 .functor NAND 1, L_0x5c7c33166ad0, L_0x5c7c33166ad0, C4<1>, C4<1>;
v0x5c7c3309ff40_0 .net "in_a", 0 0, L_0x5c7c33166ad0;  alias, 1 drivers
v0x5c7c330a0030_0 .net "in_b", 0 0, L_0x5c7c33166ad0;  alias, 1 drivers
v0x5c7c330a0120_0 .net "out", 0 0, L_0x5c7c33166b40;  alias, 1 drivers
S_0x5c7c330a07c0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c3309f0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a17f0_0 .net "in_a", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
v0x5c7c330a1890_0 .net "in_b", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
v0x5c7c330a1950_0 .net "out", 0 0, L_0x5c7c33166da0;  alias, 1 drivers
v0x5c7c330a1a70_0 .net "temp_out", 0 0, L_0x5c7c33166d30;  1 drivers
S_0x5c7c330a09a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330a07c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166d30 .functor NAND 1, L_0x5c7c33166a60, L_0x5c7c33166a60, C4<1>, C4<1>;
v0x5c7c330a0c10_0 .net "in_a", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
v0x5c7c330a0cd0_0 .net "in_b", 0 0, L_0x5c7c33166a60;  alias, 1 drivers
v0x5c7c330a0e20_0 .net "out", 0 0, L_0x5c7c33166d30;  alias, 1 drivers
S_0x5c7c330a0f20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330a07c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a1640_0 .net "in_a", 0 0, L_0x5c7c33166d30;  alias, 1 drivers
v0x5c7c330a16e0_0 .net "out", 0 0, L_0x5c7c33166da0;  alias, 1 drivers
S_0x5c7c330a10f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a0f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166da0 .functor NAND 1, L_0x5c7c33166d30, L_0x5c7c33166d30, C4<1>, C4<1>;
v0x5c7c330a1360_0 .net "in_a", 0 0, L_0x5c7c33166d30;  alias, 1 drivers
v0x5c7c330a1450_0 .net "in_b", 0 0, L_0x5c7c33166d30;  alias, 1 drivers
v0x5c7c330a1540_0 .net "out", 0 0, L_0x5c7c33166da0;  alias, 1 drivers
S_0x5c7c330a1be0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c3309f0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a2c20_0 .net "in_a", 0 0, L_0x5c7c33166bb0;  alias, 1 drivers
v0x5c7c330a2cf0_0 .net "in_b", 0 0, L_0x5c7c33166e10;  alias, 1 drivers
v0x5c7c330a2dc0_0 .net "out", 0 0, L_0x5c7c33167000;  alias, 1 drivers
v0x5c7c330a2ee0_0 .net "temp_out", 0 0, L_0x5c7c33166f90;  1 drivers
S_0x5c7c330a1dc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330a1be0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166f90 .functor NAND 1, L_0x5c7c33166bb0, L_0x5c7c33166e10, C4<1>, C4<1>;
v0x5c7c330a2010_0 .net "in_a", 0 0, L_0x5c7c33166bb0;  alias, 1 drivers
v0x5c7c330a20f0_0 .net "in_b", 0 0, L_0x5c7c33166e10;  alias, 1 drivers
v0x5c7c330a21b0_0 .net "out", 0 0, L_0x5c7c33166f90;  alias, 1 drivers
S_0x5c7c330a2300 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330a1be0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a2a70_0 .net "in_a", 0 0, L_0x5c7c33166f90;  alias, 1 drivers
v0x5c7c330a2b10_0 .net "out", 0 0, L_0x5c7c33167000;  alias, 1 drivers
S_0x5c7c330a2520 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a2300;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167000 .functor NAND 1, L_0x5c7c33166f90, L_0x5c7c33166f90, C4<1>, C4<1>;
v0x5c7c330a2790_0 .net "in_a", 0 0, L_0x5c7c33166f90;  alias, 1 drivers
v0x5c7c330a2880_0 .net "in_b", 0 0, L_0x5c7c33166f90;  alias, 1 drivers
v0x5c7c330a2970_0 .net "out", 0 0, L_0x5c7c33167000;  alias, 1 drivers
S_0x5c7c330a3030 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c3309f0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a3760_0 .net "in_a", 0 0, L_0x5c7c33166b40;  alias, 1 drivers
v0x5c7c330a3800_0 .net "out", 0 0, L_0x5c7c33166bb0;  alias, 1 drivers
S_0x5c7c330a3200 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a3030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166bb0 .functor NAND 1, L_0x5c7c33166b40, L_0x5c7c33166b40, C4<1>, C4<1>;
v0x5c7c330a3470_0 .net "in_a", 0 0, L_0x5c7c33166b40;  alias, 1 drivers
v0x5c7c330a3530_0 .net "in_b", 0 0, L_0x5c7c33166b40;  alias, 1 drivers
v0x5c7c330a3680_0 .net "out", 0 0, L_0x5c7c33166bb0;  alias, 1 drivers
S_0x5c7c330a3900 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c3309f0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a40d0_0 .net "in_a", 0 0, L_0x5c7c33166da0;  alias, 1 drivers
v0x5c7c330a4170_0 .net "out", 0 0, L_0x5c7c33166e10;  alias, 1 drivers
S_0x5c7c330a3b70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a3900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33166e10 .functor NAND 1, L_0x5c7c33166da0, L_0x5c7c33166da0, C4<1>, C4<1>;
v0x5c7c330a3de0_0 .net "in_a", 0 0, L_0x5c7c33166da0;  alias, 1 drivers
v0x5c7c330a3ea0_0 .net "in_b", 0 0, L_0x5c7c33166da0;  alias, 1 drivers
v0x5c7c330a3ff0_0 .net "out", 0 0, L_0x5c7c33166e10;  alias, 1 drivers
S_0x5c7c330a4270 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c3309f0e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a4a10_0 .net "in_a", 0 0, L_0x5c7c33167000;  alias, 1 drivers
v0x5c7c330a4ab0_0 .net "out", 0 0, L_0x5c7c33167070;  alias, 1 drivers
S_0x5c7c330a4490 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a4270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167070 .functor NAND 1, L_0x5c7c33167000, L_0x5c7c33167000, C4<1>, C4<1>;
v0x5c7c330a4700_0 .net "in_a", 0 0, L_0x5c7c33167000;  alias, 1 drivers
v0x5c7c330a47c0_0 .net "in_b", 0 0, L_0x5c7c33167000;  alias, 1 drivers
v0x5c7c330a4910_0 .net "out", 0 0, L_0x5c7c33167070;  alias, 1 drivers
S_0x5c7c330a5a50 .scope module, "mux_gate13" "Mux" 15 20, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330aedb0_0 .net "in_a", 0 0, L_0x5c7c33167f60;  1 drivers
v0x5c7c330aee50_0 .net "in_b", 0 0, L_0x5c7c33168000;  1 drivers
v0x5c7c330aef60_0 .net "out", 0 0, L_0x5c7c33167de0;  1 drivers
v0x5c7c330af000_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330af0a0_0 .net "sel_out", 0 0, L_0x5c7c33167830;  1 drivers
v0x5c7c330af220_0 .net "temp_a_out", 0 0, L_0x5c7c33167910;  1 drivers
v0x5c7c330af3d0_0 .net "temp_b_out", 0 0, L_0x5c7c331679f0;  1 drivers
S_0x5c7c330a5c50 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330a5a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a6cb0_0 .net "in_a", 0 0, L_0x5c7c33167f60;  alias, 1 drivers
v0x5c7c330a6d80_0 .net "in_b", 0 0, L_0x5c7c33167830;  alias, 1 drivers
v0x5c7c330a6e50_0 .net "out", 0 0, L_0x5c7c33167910;  alias, 1 drivers
v0x5c7c330a6f70_0 .net "temp_out", 0 0, L_0x5c7c331678a0;  1 drivers
S_0x5c7c330a5ec0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330a5c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331678a0 .functor NAND 1, L_0x5c7c33167f60, L_0x5c7c33167830, C4<1>, C4<1>;
v0x5c7c330a6130_0 .net "in_a", 0 0, L_0x5c7c33167f60;  alias, 1 drivers
v0x5c7c330a6210_0 .net "in_b", 0 0, L_0x5c7c33167830;  alias, 1 drivers
v0x5c7c330a62d0_0 .net "out", 0 0, L_0x5c7c331678a0;  alias, 1 drivers
S_0x5c7c330a63f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330a5c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a6b30_0 .net "in_a", 0 0, L_0x5c7c331678a0;  alias, 1 drivers
v0x5c7c330a6bd0_0 .net "out", 0 0, L_0x5c7c33167910;  alias, 1 drivers
S_0x5c7c330a6610 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a63f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167910 .functor NAND 1, L_0x5c7c331678a0, L_0x5c7c331678a0, C4<1>, C4<1>;
v0x5c7c330a6880_0 .net "in_a", 0 0, L_0x5c7c331678a0;  alias, 1 drivers
v0x5c7c330a6940_0 .net "in_b", 0 0, L_0x5c7c331678a0;  alias, 1 drivers
v0x5c7c330a6a30_0 .net "out", 0 0, L_0x5c7c33167910;  alias, 1 drivers
S_0x5c7c330a7030 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330a5a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a8040_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330a80e0_0 .net "in_b", 0 0, L_0x5c7c33168000;  alias, 1 drivers
v0x5c7c330a81d0_0 .net "out", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
v0x5c7c330a82f0_0 .net "temp_out", 0 0, L_0x5c7c33167980;  1 drivers
S_0x5c7c330a7210 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330a7030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167980 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33168000, C4<1>, C4<1>;
v0x5c7c330a7480_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330a7540_0 .net "in_b", 0 0, L_0x5c7c33168000;  alias, 1 drivers
v0x5c7c330a7600_0 .net "out", 0 0, L_0x5c7c33167980;  alias, 1 drivers
S_0x5c7c330a7720 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330a7030;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a7e90_0 .net "in_a", 0 0, L_0x5c7c33167980;  alias, 1 drivers
v0x5c7c330a7f30_0 .net "out", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
S_0x5c7c330a7940 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a7720;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331679f0 .functor NAND 1, L_0x5c7c33167980, L_0x5c7c33167980, C4<1>, C4<1>;
v0x5c7c330a7bb0_0 .net "in_a", 0 0, L_0x5c7c33167980;  alias, 1 drivers
v0x5c7c330a7ca0_0 .net "in_b", 0 0, L_0x5c7c33167980;  alias, 1 drivers
v0x5c7c330a7d90_0 .net "out", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
S_0x5c7c330a83b0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330a5a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a8ab0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330a8b50_0 .net "out", 0 0, L_0x5c7c33167830;  alias, 1 drivers
S_0x5c7c330a8580 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a83b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167830 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330a87d0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330a8890_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330a8950_0 .net "out", 0 0, L_0x5c7c33167830;  alias, 1 drivers
S_0x5c7c330a8c50 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330a5a50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330ae700_0 .net "branch1_out", 0 0, L_0x5c7c33167b40;  1 drivers
v0x5c7c330ae830_0 .net "branch2_out", 0 0, L_0x5c7c33167c90;  1 drivers
v0x5c7c330ae980_0 .net "in_a", 0 0, L_0x5c7c33167910;  alias, 1 drivers
v0x5c7c330aea50_0 .net "in_b", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
v0x5c7c330aeaf0_0 .net "out", 0 0, L_0x5c7c33167de0;  alias, 1 drivers
v0x5c7c330aeb90_0 .net "temp1_out", 0 0, L_0x5c7c33167ad0;  1 drivers
v0x5c7c330aec30_0 .net "temp2_out", 0 0, L_0x5c7c33167c20;  1 drivers
v0x5c7c330aecd0_0 .net "temp3_out", 0 0, L_0x5c7c33167d70;  1 drivers
S_0x5c7c330a8e80 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330a8c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330a9f40_0 .net "in_a", 0 0, L_0x5c7c33167910;  alias, 1 drivers
v0x5c7c330a9fe0_0 .net "in_b", 0 0, L_0x5c7c33167910;  alias, 1 drivers
v0x5c7c330aa0a0_0 .net "out", 0 0, L_0x5c7c33167ad0;  alias, 1 drivers
v0x5c7c330aa1c0_0 .net "temp_out", 0 0, L_0x5c7c33167a60;  1 drivers
S_0x5c7c330a90f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330a8e80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167a60 .functor NAND 1, L_0x5c7c33167910, L_0x5c7c33167910, C4<1>, C4<1>;
v0x5c7c330a9360_0 .net "in_a", 0 0, L_0x5c7c33167910;  alias, 1 drivers
v0x5c7c330a9420_0 .net "in_b", 0 0, L_0x5c7c33167910;  alias, 1 drivers
v0x5c7c330a9570_0 .net "out", 0 0, L_0x5c7c33167a60;  alias, 1 drivers
S_0x5c7c330a9670 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330a8e80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330a9d90_0 .net "in_a", 0 0, L_0x5c7c33167a60;  alias, 1 drivers
v0x5c7c330a9e30_0 .net "out", 0 0, L_0x5c7c33167ad0;  alias, 1 drivers
S_0x5c7c330a9840 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330a9670;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167ad0 .functor NAND 1, L_0x5c7c33167a60, L_0x5c7c33167a60, C4<1>, C4<1>;
v0x5c7c330a9ab0_0 .net "in_a", 0 0, L_0x5c7c33167a60;  alias, 1 drivers
v0x5c7c330a9ba0_0 .net "in_b", 0 0, L_0x5c7c33167a60;  alias, 1 drivers
v0x5c7c330a9c90_0 .net "out", 0 0, L_0x5c7c33167ad0;  alias, 1 drivers
S_0x5c7c330aa330 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330a8c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330ab360_0 .net "in_a", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
v0x5c7c330ab400_0 .net "in_b", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
v0x5c7c330ab4c0_0 .net "out", 0 0, L_0x5c7c33167c20;  alias, 1 drivers
v0x5c7c330ab5e0_0 .net "temp_out", 0 0, L_0x5c7c33167bb0;  1 drivers
S_0x5c7c330aa510 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330aa330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167bb0 .functor NAND 1, L_0x5c7c331679f0, L_0x5c7c331679f0, C4<1>, C4<1>;
v0x5c7c330aa780_0 .net "in_a", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
v0x5c7c330aa840_0 .net "in_b", 0 0, L_0x5c7c331679f0;  alias, 1 drivers
v0x5c7c330aa990_0 .net "out", 0 0, L_0x5c7c33167bb0;  alias, 1 drivers
S_0x5c7c330aaa90 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330aa330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ab1b0_0 .net "in_a", 0 0, L_0x5c7c33167bb0;  alias, 1 drivers
v0x5c7c330ab250_0 .net "out", 0 0, L_0x5c7c33167c20;  alias, 1 drivers
S_0x5c7c330aac60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330aaa90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167c20 .functor NAND 1, L_0x5c7c33167bb0, L_0x5c7c33167bb0, C4<1>, C4<1>;
v0x5c7c330aaed0_0 .net "in_a", 0 0, L_0x5c7c33167bb0;  alias, 1 drivers
v0x5c7c330aafc0_0 .net "in_b", 0 0, L_0x5c7c33167bb0;  alias, 1 drivers
v0x5c7c330ab0b0_0 .net "out", 0 0, L_0x5c7c33167c20;  alias, 1 drivers
S_0x5c7c330ab750 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330a8c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330ac790_0 .net "in_a", 0 0, L_0x5c7c33167b40;  alias, 1 drivers
v0x5c7c330ac860_0 .net "in_b", 0 0, L_0x5c7c33167c90;  alias, 1 drivers
v0x5c7c330ac930_0 .net "out", 0 0, L_0x5c7c33167d70;  alias, 1 drivers
v0x5c7c330aca50_0 .net "temp_out", 0 0, L_0x5c7c33167d00;  1 drivers
S_0x5c7c330ab930 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330ab750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167d00 .functor NAND 1, L_0x5c7c33167b40, L_0x5c7c33167c90, C4<1>, C4<1>;
v0x5c7c330abb80_0 .net "in_a", 0 0, L_0x5c7c33167b40;  alias, 1 drivers
v0x5c7c330abc60_0 .net "in_b", 0 0, L_0x5c7c33167c90;  alias, 1 drivers
v0x5c7c330abd20_0 .net "out", 0 0, L_0x5c7c33167d00;  alias, 1 drivers
S_0x5c7c330abe70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330ab750;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ac5e0_0 .net "in_a", 0 0, L_0x5c7c33167d00;  alias, 1 drivers
v0x5c7c330ac680_0 .net "out", 0 0, L_0x5c7c33167d70;  alias, 1 drivers
S_0x5c7c330ac090 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330abe70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167d70 .functor NAND 1, L_0x5c7c33167d00, L_0x5c7c33167d00, C4<1>, C4<1>;
v0x5c7c330ac300_0 .net "in_a", 0 0, L_0x5c7c33167d00;  alias, 1 drivers
v0x5c7c330ac3f0_0 .net "in_b", 0 0, L_0x5c7c33167d00;  alias, 1 drivers
v0x5c7c330ac4e0_0 .net "out", 0 0, L_0x5c7c33167d70;  alias, 1 drivers
S_0x5c7c330acba0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330a8c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ad2d0_0 .net "in_a", 0 0, L_0x5c7c33167ad0;  alias, 1 drivers
v0x5c7c330ad370_0 .net "out", 0 0, L_0x5c7c33167b40;  alias, 1 drivers
S_0x5c7c330acd70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330acba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167b40 .functor NAND 1, L_0x5c7c33167ad0, L_0x5c7c33167ad0, C4<1>, C4<1>;
v0x5c7c330acfe0_0 .net "in_a", 0 0, L_0x5c7c33167ad0;  alias, 1 drivers
v0x5c7c330ad0a0_0 .net "in_b", 0 0, L_0x5c7c33167ad0;  alias, 1 drivers
v0x5c7c330ad1f0_0 .net "out", 0 0, L_0x5c7c33167b40;  alias, 1 drivers
S_0x5c7c330ad470 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330a8c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330adc40_0 .net "in_a", 0 0, L_0x5c7c33167c20;  alias, 1 drivers
v0x5c7c330adce0_0 .net "out", 0 0, L_0x5c7c33167c90;  alias, 1 drivers
S_0x5c7c330ad6e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ad470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167c90 .functor NAND 1, L_0x5c7c33167c20, L_0x5c7c33167c20, C4<1>, C4<1>;
v0x5c7c330ad950_0 .net "in_a", 0 0, L_0x5c7c33167c20;  alias, 1 drivers
v0x5c7c330ada10_0 .net "in_b", 0 0, L_0x5c7c33167c20;  alias, 1 drivers
v0x5c7c330adb60_0 .net "out", 0 0, L_0x5c7c33167c90;  alias, 1 drivers
S_0x5c7c330adde0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330a8c50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ae580_0 .net "in_a", 0 0, L_0x5c7c33167d70;  alias, 1 drivers
v0x5c7c330ae620_0 .net "out", 0 0, L_0x5c7c33167de0;  alias, 1 drivers
S_0x5c7c330ae000 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330adde0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33167de0 .functor NAND 1, L_0x5c7c33167d70, L_0x5c7c33167d70, C4<1>, C4<1>;
v0x5c7c330ae270_0 .net "in_a", 0 0, L_0x5c7c33167d70;  alias, 1 drivers
v0x5c7c330ae330_0 .net "in_b", 0 0, L_0x5c7c33167d70;  alias, 1 drivers
v0x5c7c330ae480_0 .net "out", 0 0, L_0x5c7c33167de0;  alias, 1 drivers
S_0x5c7c330af5c0 .scope module, "mux_gate14" "Mux" 15 21, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330b8920_0 .net "in_a", 0 0, L_0x5c7c33168d80;  1 drivers
v0x5c7c330b89c0_0 .net "in_b", 0 0, L_0x5c7c33168e20;  1 drivers
v0x5c7c330b8ad0_0 .net "out", 0 0, L_0x5c7c33168bc0;  1 drivers
v0x5c7c330b8b70_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330b8c10_0 .net "sel_out", 0 0, L_0x5c7c33168190;  1 drivers
v0x5c7c330b8d90_0 .net "temp_a_out", 0 0, L_0x5c7c33168270;  1 drivers
v0x5c7c330b8f40_0 .net "temp_b_out", 0 0, L_0x5c7c33168370;  1 drivers
S_0x5c7c330af7c0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330af5c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330b0820_0 .net "in_a", 0 0, L_0x5c7c33168d80;  alias, 1 drivers
v0x5c7c330b08f0_0 .net "in_b", 0 0, L_0x5c7c33168190;  alias, 1 drivers
v0x5c7c330b09c0_0 .net "out", 0 0, L_0x5c7c33168270;  alias, 1 drivers
v0x5c7c330b0ae0_0 .net "temp_out", 0 0, L_0x5c7c33168200;  1 drivers
S_0x5c7c330afa30 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330af7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168200 .functor NAND 1, L_0x5c7c33168d80, L_0x5c7c33168190, C4<1>, C4<1>;
v0x5c7c330afca0_0 .net "in_a", 0 0, L_0x5c7c33168d80;  alias, 1 drivers
v0x5c7c330afd80_0 .net "in_b", 0 0, L_0x5c7c33168190;  alias, 1 drivers
v0x5c7c330afe40_0 .net "out", 0 0, L_0x5c7c33168200;  alias, 1 drivers
S_0x5c7c330aff60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330af7c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b06a0_0 .net "in_a", 0 0, L_0x5c7c33168200;  alias, 1 drivers
v0x5c7c330b0740_0 .net "out", 0 0, L_0x5c7c33168270;  alias, 1 drivers
S_0x5c7c330b0180 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330aff60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168270 .functor NAND 1, L_0x5c7c33168200, L_0x5c7c33168200, C4<1>, C4<1>;
v0x5c7c330b03f0_0 .net "in_a", 0 0, L_0x5c7c33168200;  alias, 1 drivers
v0x5c7c330b04b0_0 .net "in_b", 0 0, L_0x5c7c33168200;  alias, 1 drivers
v0x5c7c330b05a0_0 .net "out", 0 0, L_0x5c7c33168270;  alias, 1 drivers
S_0x5c7c330b0ba0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330af5c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330b1bb0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330b1c50_0 .net "in_b", 0 0, L_0x5c7c33168e20;  alias, 1 drivers
v0x5c7c330b1d40_0 .net "out", 0 0, L_0x5c7c33168370;  alias, 1 drivers
v0x5c7c330b1e60_0 .net "temp_out", 0 0, L_0x5c7c331682e0;  1 drivers
S_0x5c7c330b0d80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330b0ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331682e0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33168e20, C4<1>, C4<1>;
v0x5c7c330b0ff0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330b10b0_0 .net "in_b", 0 0, L_0x5c7c33168e20;  alias, 1 drivers
v0x5c7c330b1170_0 .net "out", 0 0, L_0x5c7c331682e0;  alias, 1 drivers
S_0x5c7c330b1290 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330b0ba0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b1a00_0 .net "in_a", 0 0, L_0x5c7c331682e0;  alias, 1 drivers
v0x5c7c330b1aa0_0 .net "out", 0 0, L_0x5c7c33168370;  alias, 1 drivers
S_0x5c7c330b14b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b1290;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168370 .functor NAND 1, L_0x5c7c331682e0, L_0x5c7c331682e0, C4<1>, C4<1>;
v0x5c7c330b1720_0 .net "in_a", 0 0, L_0x5c7c331682e0;  alias, 1 drivers
v0x5c7c330b1810_0 .net "in_b", 0 0, L_0x5c7c331682e0;  alias, 1 drivers
v0x5c7c330b1900_0 .net "out", 0 0, L_0x5c7c33168370;  alias, 1 drivers
S_0x5c7c330b1f20 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330af5c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b2620_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330b26c0_0 .net "out", 0 0, L_0x5c7c33168190;  alias, 1 drivers
S_0x5c7c330b20f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b1f20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168190 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330b2340_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330b2400_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330b24c0_0 .net "out", 0 0, L_0x5c7c33168190;  alias, 1 drivers
S_0x5c7c330b27c0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330af5c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330b8270_0 .net "branch1_out", 0 0, L_0x5c7c33168580;  1 drivers
v0x5c7c330b83a0_0 .net "branch2_out", 0 0, L_0x5c7c331688a0;  1 drivers
v0x5c7c330b84f0_0 .net "in_a", 0 0, L_0x5c7c33168270;  alias, 1 drivers
v0x5c7c330b85c0_0 .net "in_b", 0 0, L_0x5c7c33168370;  alias, 1 drivers
v0x5c7c330b8660_0 .net "out", 0 0, L_0x5c7c33168bc0;  alias, 1 drivers
v0x5c7c330b8700_0 .net "temp1_out", 0 0, L_0x5c7c331684d0;  1 drivers
v0x5c7c330b87a0_0 .net "temp2_out", 0 0, L_0x5c7c331687f0;  1 drivers
v0x5c7c330b8840_0 .net "temp3_out", 0 0, L_0x5c7c33168b10;  1 drivers
S_0x5c7c330b29f0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330b27c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330b3ab0_0 .net "in_a", 0 0, L_0x5c7c33168270;  alias, 1 drivers
v0x5c7c330b3b50_0 .net "in_b", 0 0, L_0x5c7c33168270;  alias, 1 drivers
v0x5c7c330b3c10_0 .net "out", 0 0, L_0x5c7c331684d0;  alias, 1 drivers
v0x5c7c330b3d30_0 .net "temp_out", 0 0, L_0x5c7c33168420;  1 drivers
S_0x5c7c330b2c60 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330b29f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168420 .functor NAND 1, L_0x5c7c33168270, L_0x5c7c33168270, C4<1>, C4<1>;
v0x5c7c330b2ed0_0 .net "in_a", 0 0, L_0x5c7c33168270;  alias, 1 drivers
v0x5c7c330b2f90_0 .net "in_b", 0 0, L_0x5c7c33168270;  alias, 1 drivers
v0x5c7c330b30e0_0 .net "out", 0 0, L_0x5c7c33168420;  alias, 1 drivers
S_0x5c7c330b31e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330b29f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b3900_0 .net "in_a", 0 0, L_0x5c7c33168420;  alias, 1 drivers
v0x5c7c330b39a0_0 .net "out", 0 0, L_0x5c7c331684d0;  alias, 1 drivers
S_0x5c7c330b33b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b31e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331684d0 .functor NAND 1, L_0x5c7c33168420, L_0x5c7c33168420, C4<1>, C4<1>;
v0x5c7c330b3620_0 .net "in_a", 0 0, L_0x5c7c33168420;  alias, 1 drivers
v0x5c7c330b3710_0 .net "in_b", 0 0, L_0x5c7c33168420;  alias, 1 drivers
v0x5c7c330b3800_0 .net "out", 0 0, L_0x5c7c331684d0;  alias, 1 drivers
S_0x5c7c330b3ea0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330b27c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330b4ed0_0 .net "in_a", 0 0, L_0x5c7c33168370;  alias, 1 drivers
v0x5c7c330b4f70_0 .net "in_b", 0 0, L_0x5c7c33168370;  alias, 1 drivers
v0x5c7c330b5030_0 .net "out", 0 0, L_0x5c7c331687f0;  alias, 1 drivers
v0x5c7c330b5150_0 .net "temp_out", 0 0, L_0x5c7c33168740;  1 drivers
S_0x5c7c330b4080 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330b3ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168740 .functor NAND 1, L_0x5c7c33168370, L_0x5c7c33168370, C4<1>, C4<1>;
v0x5c7c330b42f0_0 .net "in_a", 0 0, L_0x5c7c33168370;  alias, 1 drivers
v0x5c7c330b43b0_0 .net "in_b", 0 0, L_0x5c7c33168370;  alias, 1 drivers
v0x5c7c330b4500_0 .net "out", 0 0, L_0x5c7c33168740;  alias, 1 drivers
S_0x5c7c330b4600 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330b3ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b4d20_0 .net "in_a", 0 0, L_0x5c7c33168740;  alias, 1 drivers
v0x5c7c330b4dc0_0 .net "out", 0 0, L_0x5c7c331687f0;  alias, 1 drivers
S_0x5c7c330b47d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b4600;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331687f0 .functor NAND 1, L_0x5c7c33168740, L_0x5c7c33168740, C4<1>, C4<1>;
v0x5c7c330b4a40_0 .net "in_a", 0 0, L_0x5c7c33168740;  alias, 1 drivers
v0x5c7c330b4b30_0 .net "in_b", 0 0, L_0x5c7c33168740;  alias, 1 drivers
v0x5c7c330b4c20_0 .net "out", 0 0, L_0x5c7c331687f0;  alias, 1 drivers
S_0x5c7c330b52c0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330b27c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330b6300_0 .net "in_a", 0 0, L_0x5c7c33168580;  alias, 1 drivers
v0x5c7c330b63d0_0 .net "in_b", 0 0, L_0x5c7c331688a0;  alias, 1 drivers
v0x5c7c330b64a0_0 .net "out", 0 0, L_0x5c7c33168b10;  alias, 1 drivers
v0x5c7c330b65c0_0 .net "temp_out", 0 0, L_0x5c7c33168a60;  1 drivers
S_0x5c7c330b54a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330b52c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168a60 .functor NAND 1, L_0x5c7c33168580, L_0x5c7c331688a0, C4<1>, C4<1>;
v0x5c7c330b56f0_0 .net "in_a", 0 0, L_0x5c7c33168580;  alias, 1 drivers
v0x5c7c330b57d0_0 .net "in_b", 0 0, L_0x5c7c331688a0;  alias, 1 drivers
v0x5c7c330b5890_0 .net "out", 0 0, L_0x5c7c33168a60;  alias, 1 drivers
S_0x5c7c330b59e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330b52c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b6150_0 .net "in_a", 0 0, L_0x5c7c33168a60;  alias, 1 drivers
v0x5c7c330b61f0_0 .net "out", 0 0, L_0x5c7c33168b10;  alias, 1 drivers
S_0x5c7c330b5c00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b59e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168b10 .functor NAND 1, L_0x5c7c33168a60, L_0x5c7c33168a60, C4<1>, C4<1>;
v0x5c7c330b5e70_0 .net "in_a", 0 0, L_0x5c7c33168a60;  alias, 1 drivers
v0x5c7c330b5f60_0 .net "in_b", 0 0, L_0x5c7c33168a60;  alias, 1 drivers
v0x5c7c330b6050_0 .net "out", 0 0, L_0x5c7c33168b10;  alias, 1 drivers
S_0x5c7c330b6710 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330b27c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b6e40_0 .net "in_a", 0 0, L_0x5c7c331684d0;  alias, 1 drivers
v0x5c7c330b6ee0_0 .net "out", 0 0, L_0x5c7c33168580;  alias, 1 drivers
S_0x5c7c330b68e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b6710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168580 .functor NAND 1, L_0x5c7c331684d0, L_0x5c7c331684d0, C4<1>, C4<1>;
v0x5c7c330b6b50_0 .net "in_a", 0 0, L_0x5c7c331684d0;  alias, 1 drivers
v0x5c7c330b6c10_0 .net "in_b", 0 0, L_0x5c7c331684d0;  alias, 1 drivers
v0x5c7c330b6d60_0 .net "out", 0 0, L_0x5c7c33168580;  alias, 1 drivers
S_0x5c7c330b6fe0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330b27c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b77b0_0 .net "in_a", 0 0, L_0x5c7c331687f0;  alias, 1 drivers
v0x5c7c330b7850_0 .net "out", 0 0, L_0x5c7c331688a0;  alias, 1 drivers
S_0x5c7c330b7250 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b6fe0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331688a0 .functor NAND 1, L_0x5c7c331687f0, L_0x5c7c331687f0, C4<1>, C4<1>;
v0x5c7c330b74c0_0 .net "in_a", 0 0, L_0x5c7c331687f0;  alias, 1 drivers
v0x5c7c330b7580_0 .net "in_b", 0 0, L_0x5c7c331687f0;  alias, 1 drivers
v0x5c7c330b76d0_0 .net "out", 0 0, L_0x5c7c331688a0;  alias, 1 drivers
S_0x5c7c330b7950 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330b27c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330b80f0_0 .net "in_a", 0 0, L_0x5c7c33168b10;  alias, 1 drivers
v0x5c7c330b8190_0 .net "out", 0 0, L_0x5c7c33168bc0;  alias, 1 drivers
S_0x5c7c330b7b70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b7950;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168bc0 .functor NAND 1, L_0x5c7c33168b10, L_0x5c7c33168b10, C4<1>, C4<1>;
v0x5c7c330b7de0_0 .net "in_a", 0 0, L_0x5c7c33168b10;  alias, 1 drivers
v0x5c7c330b7ea0_0 .net "in_b", 0 0, L_0x5c7c33168b10;  alias, 1 drivers
v0x5c7c330b7ff0_0 .net "out", 0 0, L_0x5c7c33168bc0;  alias, 1 drivers
S_0x5c7c330b9130 .scope module, "mux_gate15" "Mux" 15 22, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330c2490_0 .net "in_a", 0 0, L_0x5c7c33169c90;  1 drivers
v0x5c7c330c2530_0 .net "in_b", 0 0, L_0x5c7c33169d30;  1 drivers
v0x5c7c330c2640_0 .net "out", 0 0, L_0x5c7c33169ad0;  1 drivers
v0x5c7c330c26e0_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330c2780_0 .net "sel_out", 0 0, L_0x5c7c33168fc0;  1 drivers
v0x5c7c330c2900_0 .net "temp_a_out", 0 0, L_0x5c7c33169120;  1 drivers
v0x5c7c330c2ab0_0 .net "temp_b_out", 0 0, L_0x5c7c33169280;  1 drivers
S_0x5c7c330b9330 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330b9130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330ba390_0 .net "in_a", 0 0, L_0x5c7c33169c90;  alias, 1 drivers
v0x5c7c330ba460_0 .net "in_b", 0 0, L_0x5c7c33168fc0;  alias, 1 drivers
v0x5c7c330ba530_0 .net "out", 0 0, L_0x5c7c33169120;  alias, 1 drivers
v0x5c7c330ba650_0 .net "temp_out", 0 0, L_0x5c7c33169070;  1 drivers
S_0x5c7c330b95a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330b9330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169070 .functor NAND 1, L_0x5c7c33169c90, L_0x5c7c33168fc0, C4<1>, C4<1>;
v0x5c7c330b9810_0 .net "in_a", 0 0, L_0x5c7c33169c90;  alias, 1 drivers
v0x5c7c330b98f0_0 .net "in_b", 0 0, L_0x5c7c33168fc0;  alias, 1 drivers
v0x5c7c330b99b0_0 .net "out", 0 0, L_0x5c7c33169070;  alias, 1 drivers
S_0x5c7c330b9ad0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330b9330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ba210_0 .net "in_a", 0 0, L_0x5c7c33169070;  alias, 1 drivers
v0x5c7c330ba2b0_0 .net "out", 0 0, L_0x5c7c33169120;  alias, 1 drivers
S_0x5c7c330b9cf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330b9ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169120 .functor NAND 1, L_0x5c7c33169070, L_0x5c7c33169070, C4<1>, C4<1>;
v0x5c7c330b9f60_0 .net "in_a", 0 0, L_0x5c7c33169070;  alias, 1 drivers
v0x5c7c330ba020_0 .net "in_b", 0 0, L_0x5c7c33169070;  alias, 1 drivers
v0x5c7c330ba110_0 .net "out", 0 0, L_0x5c7c33169120;  alias, 1 drivers
S_0x5c7c330ba710 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330b9130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330bb720_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330bb7c0_0 .net "in_b", 0 0, L_0x5c7c33169d30;  alias, 1 drivers
v0x5c7c330bb8b0_0 .net "out", 0 0, L_0x5c7c33169280;  alias, 1 drivers
v0x5c7c330bb9d0_0 .net "temp_out", 0 0, L_0x5c7c331691d0;  1 drivers
S_0x5c7c330ba8f0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330ba710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331691d0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169d30, C4<1>, C4<1>;
v0x5c7c330bab60_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330bac20_0 .net "in_b", 0 0, L_0x5c7c33169d30;  alias, 1 drivers
v0x5c7c330bace0_0 .net "out", 0 0, L_0x5c7c331691d0;  alias, 1 drivers
S_0x5c7c330bae00 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330ba710;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330bb570_0 .net "in_a", 0 0, L_0x5c7c331691d0;  alias, 1 drivers
v0x5c7c330bb610_0 .net "out", 0 0, L_0x5c7c33169280;  alias, 1 drivers
S_0x5c7c330bb020 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330bae00;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169280 .functor NAND 1, L_0x5c7c331691d0, L_0x5c7c331691d0, C4<1>, C4<1>;
v0x5c7c330bb290_0 .net "in_a", 0 0, L_0x5c7c331691d0;  alias, 1 drivers
v0x5c7c330bb380_0 .net "in_b", 0 0, L_0x5c7c331691d0;  alias, 1 drivers
v0x5c7c330bb470_0 .net "out", 0 0, L_0x5c7c33169280;  alias, 1 drivers
S_0x5c7c330bba90 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330b9130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330bc190_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330bc230_0 .net "out", 0 0, L_0x5c7c33168fc0;  alias, 1 drivers
S_0x5c7c330bbc60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330bba90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33168fc0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330bbeb0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330bbf70_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330bc030_0 .net "out", 0 0, L_0x5c7c33168fc0;  alias, 1 drivers
S_0x5c7c330bc330 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330b9130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330c1de0_0 .net "branch1_out", 0 0, L_0x5c7c33169490;  1 drivers
v0x5c7c330c1f10_0 .net "branch2_out", 0 0, L_0x5c7c331697b0;  1 drivers
v0x5c7c330c2060_0 .net "in_a", 0 0, L_0x5c7c33169120;  alias, 1 drivers
v0x5c7c330c2130_0 .net "in_b", 0 0, L_0x5c7c33169280;  alias, 1 drivers
v0x5c7c330c21d0_0 .net "out", 0 0, L_0x5c7c33169ad0;  alias, 1 drivers
v0x5c7c330c2270_0 .net "temp1_out", 0 0, L_0x5c7c331693e0;  1 drivers
v0x5c7c330c2310_0 .net "temp2_out", 0 0, L_0x5c7c33169700;  1 drivers
v0x5c7c330c23b0_0 .net "temp3_out", 0 0, L_0x5c7c33169a20;  1 drivers
S_0x5c7c330bc560 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330bc330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330bd620_0 .net "in_a", 0 0, L_0x5c7c33169120;  alias, 1 drivers
v0x5c7c330bd6c0_0 .net "in_b", 0 0, L_0x5c7c33169120;  alias, 1 drivers
v0x5c7c330bd780_0 .net "out", 0 0, L_0x5c7c331693e0;  alias, 1 drivers
v0x5c7c330bd8a0_0 .net "temp_out", 0 0, L_0x5c7c33169330;  1 drivers
S_0x5c7c330bc7d0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330bc560;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169330 .functor NAND 1, L_0x5c7c33169120, L_0x5c7c33169120, C4<1>, C4<1>;
v0x5c7c330bca40_0 .net "in_a", 0 0, L_0x5c7c33169120;  alias, 1 drivers
v0x5c7c330bcb00_0 .net "in_b", 0 0, L_0x5c7c33169120;  alias, 1 drivers
v0x5c7c330bcc50_0 .net "out", 0 0, L_0x5c7c33169330;  alias, 1 drivers
S_0x5c7c330bcd50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330bc560;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330bd470_0 .net "in_a", 0 0, L_0x5c7c33169330;  alias, 1 drivers
v0x5c7c330bd510_0 .net "out", 0 0, L_0x5c7c331693e0;  alias, 1 drivers
S_0x5c7c330bcf20 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330bcd50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331693e0 .functor NAND 1, L_0x5c7c33169330, L_0x5c7c33169330, C4<1>, C4<1>;
v0x5c7c330bd190_0 .net "in_a", 0 0, L_0x5c7c33169330;  alias, 1 drivers
v0x5c7c330bd280_0 .net "in_b", 0 0, L_0x5c7c33169330;  alias, 1 drivers
v0x5c7c330bd370_0 .net "out", 0 0, L_0x5c7c331693e0;  alias, 1 drivers
S_0x5c7c330bda10 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330bc330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330bea40_0 .net "in_a", 0 0, L_0x5c7c33169280;  alias, 1 drivers
v0x5c7c330beae0_0 .net "in_b", 0 0, L_0x5c7c33169280;  alias, 1 drivers
v0x5c7c330beba0_0 .net "out", 0 0, L_0x5c7c33169700;  alias, 1 drivers
v0x5c7c330becc0_0 .net "temp_out", 0 0, L_0x5c7c33169650;  1 drivers
S_0x5c7c330bdbf0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330bda10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169650 .functor NAND 1, L_0x5c7c33169280, L_0x5c7c33169280, C4<1>, C4<1>;
v0x5c7c330bde60_0 .net "in_a", 0 0, L_0x5c7c33169280;  alias, 1 drivers
v0x5c7c330bdf20_0 .net "in_b", 0 0, L_0x5c7c33169280;  alias, 1 drivers
v0x5c7c330be070_0 .net "out", 0 0, L_0x5c7c33169650;  alias, 1 drivers
S_0x5c7c330be170 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330bda10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330be890_0 .net "in_a", 0 0, L_0x5c7c33169650;  alias, 1 drivers
v0x5c7c330be930_0 .net "out", 0 0, L_0x5c7c33169700;  alias, 1 drivers
S_0x5c7c330be340 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330be170;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169700 .functor NAND 1, L_0x5c7c33169650, L_0x5c7c33169650, C4<1>, C4<1>;
v0x5c7c330be5b0_0 .net "in_a", 0 0, L_0x5c7c33169650;  alias, 1 drivers
v0x5c7c330be6a0_0 .net "in_b", 0 0, L_0x5c7c33169650;  alias, 1 drivers
v0x5c7c330be790_0 .net "out", 0 0, L_0x5c7c33169700;  alias, 1 drivers
S_0x5c7c330bee30 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330bc330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330bfe70_0 .net "in_a", 0 0, L_0x5c7c33169490;  alias, 1 drivers
v0x5c7c330bff40_0 .net "in_b", 0 0, L_0x5c7c331697b0;  alias, 1 drivers
v0x5c7c330c0010_0 .net "out", 0 0, L_0x5c7c33169a20;  alias, 1 drivers
v0x5c7c330c0130_0 .net "temp_out", 0 0, L_0x5c7c33169970;  1 drivers
S_0x5c7c330bf010 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330bee30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169970 .functor NAND 1, L_0x5c7c33169490, L_0x5c7c331697b0, C4<1>, C4<1>;
v0x5c7c330bf260_0 .net "in_a", 0 0, L_0x5c7c33169490;  alias, 1 drivers
v0x5c7c330bf340_0 .net "in_b", 0 0, L_0x5c7c331697b0;  alias, 1 drivers
v0x5c7c330bf400_0 .net "out", 0 0, L_0x5c7c33169970;  alias, 1 drivers
S_0x5c7c330bf550 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330bee30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330bfcc0_0 .net "in_a", 0 0, L_0x5c7c33169970;  alias, 1 drivers
v0x5c7c330bfd60_0 .net "out", 0 0, L_0x5c7c33169a20;  alias, 1 drivers
S_0x5c7c330bf770 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330bf550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169a20 .functor NAND 1, L_0x5c7c33169970, L_0x5c7c33169970, C4<1>, C4<1>;
v0x5c7c330bf9e0_0 .net "in_a", 0 0, L_0x5c7c33169970;  alias, 1 drivers
v0x5c7c330bfad0_0 .net "in_b", 0 0, L_0x5c7c33169970;  alias, 1 drivers
v0x5c7c330bfbc0_0 .net "out", 0 0, L_0x5c7c33169a20;  alias, 1 drivers
S_0x5c7c330c0280 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330bc330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c09b0_0 .net "in_a", 0 0, L_0x5c7c331693e0;  alias, 1 drivers
v0x5c7c330c0a50_0 .net "out", 0 0, L_0x5c7c33169490;  alias, 1 drivers
S_0x5c7c330c0450 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c0280;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169490 .functor NAND 1, L_0x5c7c331693e0, L_0x5c7c331693e0, C4<1>, C4<1>;
v0x5c7c330c06c0_0 .net "in_a", 0 0, L_0x5c7c331693e0;  alias, 1 drivers
v0x5c7c330c0780_0 .net "in_b", 0 0, L_0x5c7c331693e0;  alias, 1 drivers
v0x5c7c330c08d0_0 .net "out", 0 0, L_0x5c7c33169490;  alias, 1 drivers
S_0x5c7c330c0b50 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330bc330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c1320_0 .net "in_a", 0 0, L_0x5c7c33169700;  alias, 1 drivers
v0x5c7c330c13c0_0 .net "out", 0 0, L_0x5c7c331697b0;  alias, 1 drivers
S_0x5c7c330c0dc0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c0b50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331697b0 .functor NAND 1, L_0x5c7c33169700, L_0x5c7c33169700, C4<1>, C4<1>;
v0x5c7c330c1030_0 .net "in_a", 0 0, L_0x5c7c33169700;  alias, 1 drivers
v0x5c7c330c10f0_0 .net "in_b", 0 0, L_0x5c7c33169700;  alias, 1 drivers
v0x5c7c330c1240_0 .net "out", 0 0, L_0x5c7c331697b0;  alias, 1 drivers
S_0x5c7c330c14c0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330bc330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c1c60_0 .net "in_a", 0 0, L_0x5c7c33169a20;  alias, 1 drivers
v0x5c7c330c1d00_0 .net "out", 0 0, L_0x5c7c33169ad0;  alias, 1 drivers
S_0x5c7c330c16e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c14c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33169ad0 .functor NAND 1, L_0x5c7c33169a20, L_0x5c7c33169a20, C4<1>, C4<1>;
v0x5c7c330c1950_0 .net "in_a", 0 0, L_0x5c7c33169a20;  alias, 1 drivers
v0x5c7c330c1a10_0 .net "in_b", 0 0, L_0x5c7c33169a20;  alias, 1 drivers
v0x5c7c330c1b60_0 .net "out", 0 0, L_0x5c7c33169ad0;  alias, 1 drivers
S_0x5c7c330c2ca0 .scope module, "mux_gate2" "Mux" 15 9, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330cc040_0 .net "in_a", 0 0, L_0x5c7c3315df00;  1 drivers
v0x5c7c330cc0e0_0 .net "in_b", 0 0, L_0x5c7c3315dfa0;  1 drivers
v0x5c7c330cc1f0_0 .net "out", 0 0, L_0x5c7c3315dd40;  1 drivers
v0x5c7c330cc290_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330cc330_0 .net "sel_out", 0 0, L_0x5c7c3315d250;  1 drivers
v0x5c7c330cc4b0_0 .net "temp_a_out", 0 0, L_0x5c7c3315d390;  1 drivers
v0x5c7c330cc660_0 .net "temp_b_out", 0 0, L_0x5c7c3315d4f0;  1 drivers
S_0x5c7c330c2ea0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330c2ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330c3eb0_0 .net "in_a", 0 0, L_0x5c7c3315df00;  alias, 1 drivers
v0x5c7c330c3f80_0 .net "in_b", 0 0, L_0x5c7c3315d250;  alias, 1 drivers
v0x5c7c330c4050_0 .net "out", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
v0x5c7c330c4170_0 .net "temp_out", 0 0, L_0x5c7c3315d2e0;  1 drivers
S_0x5c7c330c30c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330c2ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d2e0 .functor NAND 1, L_0x5c7c3315df00, L_0x5c7c3315d250, C4<1>, C4<1>;
v0x5c7c330c3330_0 .net "in_a", 0 0, L_0x5c7c3315df00;  alias, 1 drivers
v0x5c7c330c3410_0 .net "in_b", 0 0, L_0x5c7c3315d250;  alias, 1 drivers
v0x5c7c330c34d0_0 .net "out", 0 0, L_0x5c7c3315d2e0;  alias, 1 drivers
S_0x5c7c330c35f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330c2ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c3d30_0 .net "in_a", 0 0, L_0x5c7c3315d2e0;  alias, 1 drivers
v0x5c7c330c3dd0_0 .net "out", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
S_0x5c7c330c3810 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c35f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d390 .functor NAND 1, L_0x5c7c3315d2e0, L_0x5c7c3315d2e0, C4<1>, C4<1>;
v0x5c7c330c3a80_0 .net "in_a", 0 0, L_0x5c7c3315d2e0;  alias, 1 drivers
v0x5c7c330c3b40_0 .net "in_b", 0 0, L_0x5c7c3315d2e0;  alias, 1 drivers
v0x5c7c330c3c30_0 .net "out", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
S_0x5c7c330c4230 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330c2ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330c5240_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330c52e0_0 .net "in_b", 0 0, L_0x5c7c3315dfa0;  alias, 1 drivers
v0x5c7c330c53d0_0 .net "out", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
v0x5c7c330c54f0_0 .net "temp_out", 0 0, L_0x5c7c3315d440;  1 drivers
S_0x5c7c330c4410 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330c4230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d440 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c3315dfa0, C4<1>, C4<1>;
v0x5c7c330c4680_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330c4740_0 .net "in_b", 0 0, L_0x5c7c3315dfa0;  alias, 1 drivers
v0x5c7c330c4800_0 .net "out", 0 0, L_0x5c7c3315d440;  alias, 1 drivers
S_0x5c7c330c4920 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330c4230;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c5090_0 .net "in_a", 0 0, L_0x5c7c3315d440;  alias, 1 drivers
v0x5c7c330c5130_0 .net "out", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
S_0x5c7c330c4b40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c4920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d4f0 .functor NAND 1, L_0x5c7c3315d440, L_0x5c7c3315d440, C4<1>, C4<1>;
v0x5c7c330c4db0_0 .net "in_a", 0 0, L_0x5c7c3315d440;  alias, 1 drivers
v0x5c7c330c4ea0_0 .net "in_b", 0 0, L_0x5c7c3315d440;  alias, 1 drivers
v0x5c7c330c4f90_0 .net "out", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
S_0x5c7c330c5640 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330c2ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c5d40_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330c5de0_0 .net "out", 0 0, L_0x5c7c3315d250;  alias, 1 drivers
S_0x5c7c330c5810 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c5640;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d250 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330c5a60_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330c5b20_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330c5be0_0 .net "out", 0 0, L_0x5c7c3315d250;  alias, 1 drivers
S_0x5c7c330c5ee0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330c2ca0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330cb990_0 .net "branch1_out", 0 0, L_0x5c7c3315d700;  1 drivers
v0x5c7c330cbac0_0 .net "branch2_out", 0 0, L_0x5c7c3315da20;  1 drivers
v0x5c7c330cbc10_0 .net "in_a", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
v0x5c7c330cbce0_0 .net "in_b", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
v0x5c7c330cbd80_0 .net "out", 0 0, L_0x5c7c3315dd40;  alias, 1 drivers
v0x5c7c330cbe20_0 .net "temp1_out", 0 0, L_0x5c7c3315d650;  1 drivers
v0x5c7c330cbec0_0 .net "temp2_out", 0 0, L_0x5c7c3315d970;  1 drivers
v0x5c7c330cbf60_0 .net "temp3_out", 0 0, L_0x5c7c3315dc90;  1 drivers
S_0x5c7c330c6110 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330c5ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330c71d0_0 .net "in_a", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
v0x5c7c330c7270_0 .net "in_b", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
v0x5c7c330c7330_0 .net "out", 0 0, L_0x5c7c3315d650;  alias, 1 drivers
v0x5c7c330c7450_0 .net "temp_out", 0 0, L_0x5c7c3315d5a0;  1 drivers
S_0x5c7c330c6380 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330c6110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d5a0 .functor NAND 1, L_0x5c7c3315d390, L_0x5c7c3315d390, C4<1>, C4<1>;
v0x5c7c330c65f0_0 .net "in_a", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
v0x5c7c330c66b0_0 .net "in_b", 0 0, L_0x5c7c3315d390;  alias, 1 drivers
v0x5c7c330c6800_0 .net "out", 0 0, L_0x5c7c3315d5a0;  alias, 1 drivers
S_0x5c7c330c6900 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330c6110;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c7020_0 .net "in_a", 0 0, L_0x5c7c3315d5a0;  alias, 1 drivers
v0x5c7c330c70c0_0 .net "out", 0 0, L_0x5c7c3315d650;  alias, 1 drivers
S_0x5c7c330c6ad0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c6900;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d650 .functor NAND 1, L_0x5c7c3315d5a0, L_0x5c7c3315d5a0, C4<1>, C4<1>;
v0x5c7c330c6d40_0 .net "in_a", 0 0, L_0x5c7c3315d5a0;  alias, 1 drivers
v0x5c7c330c6e30_0 .net "in_b", 0 0, L_0x5c7c3315d5a0;  alias, 1 drivers
v0x5c7c330c6f20_0 .net "out", 0 0, L_0x5c7c3315d650;  alias, 1 drivers
S_0x5c7c330c75c0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330c5ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330c85f0_0 .net "in_a", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
v0x5c7c330c8690_0 .net "in_b", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
v0x5c7c330c8750_0 .net "out", 0 0, L_0x5c7c3315d970;  alias, 1 drivers
v0x5c7c330c8870_0 .net "temp_out", 0 0, L_0x5c7c3315d8c0;  1 drivers
S_0x5c7c330c77a0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330c75c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d8c0 .functor NAND 1, L_0x5c7c3315d4f0, L_0x5c7c3315d4f0, C4<1>, C4<1>;
v0x5c7c330c7a10_0 .net "in_a", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
v0x5c7c330c7ad0_0 .net "in_b", 0 0, L_0x5c7c3315d4f0;  alias, 1 drivers
v0x5c7c330c7c20_0 .net "out", 0 0, L_0x5c7c3315d8c0;  alias, 1 drivers
S_0x5c7c330c7d20 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330c75c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c8440_0 .net "in_a", 0 0, L_0x5c7c3315d8c0;  alias, 1 drivers
v0x5c7c330c84e0_0 .net "out", 0 0, L_0x5c7c3315d970;  alias, 1 drivers
S_0x5c7c330c7ef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c7d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d970 .functor NAND 1, L_0x5c7c3315d8c0, L_0x5c7c3315d8c0, C4<1>, C4<1>;
v0x5c7c330c8160_0 .net "in_a", 0 0, L_0x5c7c3315d8c0;  alias, 1 drivers
v0x5c7c330c8250_0 .net "in_b", 0 0, L_0x5c7c3315d8c0;  alias, 1 drivers
v0x5c7c330c8340_0 .net "out", 0 0, L_0x5c7c3315d970;  alias, 1 drivers
S_0x5c7c330c89e0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330c5ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330c9a20_0 .net "in_a", 0 0, L_0x5c7c3315d700;  alias, 1 drivers
v0x5c7c330c9af0_0 .net "in_b", 0 0, L_0x5c7c3315da20;  alias, 1 drivers
v0x5c7c330c9bc0_0 .net "out", 0 0, L_0x5c7c3315dc90;  alias, 1 drivers
v0x5c7c330c9ce0_0 .net "temp_out", 0 0, L_0x5c7c3315dbe0;  1 drivers
S_0x5c7c330c8bc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330c89e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315dbe0 .functor NAND 1, L_0x5c7c3315d700, L_0x5c7c3315da20, C4<1>, C4<1>;
v0x5c7c330c8e10_0 .net "in_a", 0 0, L_0x5c7c3315d700;  alias, 1 drivers
v0x5c7c330c8ef0_0 .net "in_b", 0 0, L_0x5c7c3315da20;  alias, 1 drivers
v0x5c7c330c8fb0_0 .net "out", 0 0, L_0x5c7c3315dbe0;  alias, 1 drivers
S_0x5c7c330c9100 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330c89e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330c9870_0 .net "in_a", 0 0, L_0x5c7c3315dbe0;  alias, 1 drivers
v0x5c7c330c9910_0 .net "out", 0 0, L_0x5c7c3315dc90;  alias, 1 drivers
S_0x5c7c330c9320 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c9100;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315dc90 .functor NAND 1, L_0x5c7c3315dbe0, L_0x5c7c3315dbe0, C4<1>, C4<1>;
v0x5c7c330c9590_0 .net "in_a", 0 0, L_0x5c7c3315dbe0;  alias, 1 drivers
v0x5c7c330c9680_0 .net "in_b", 0 0, L_0x5c7c3315dbe0;  alias, 1 drivers
v0x5c7c330c9770_0 .net "out", 0 0, L_0x5c7c3315dc90;  alias, 1 drivers
S_0x5c7c330c9e30 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330c5ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ca560_0 .net "in_a", 0 0, L_0x5c7c3315d650;  alias, 1 drivers
v0x5c7c330ca600_0 .net "out", 0 0, L_0x5c7c3315d700;  alias, 1 drivers
S_0x5c7c330ca000 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330c9e30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315d700 .functor NAND 1, L_0x5c7c3315d650, L_0x5c7c3315d650, C4<1>, C4<1>;
v0x5c7c330ca270_0 .net "in_a", 0 0, L_0x5c7c3315d650;  alias, 1 drivers
v0x5c7c330ca330_0 .net "in_b", 0 0, L_0x5c7c3315d650;  alias, 1 drivers
v0x5c7c330ca480_0 .net "out", 0 0, L_0x5c7c3315d700;  alias, 1 drivers
S_0x5c7c330ca700 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330c5ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330caed0_0 .net "in_a", 0 0, L_0x5c7c3315d970;  alias, 1 drivers
v0x5c7c330caf70_0 .net "out", 0 0, L_0x5c7c3315da20;  alias, 1 drivers
S_0x5c7c330ca970 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ca700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315da20 .functor NAND 1, L_0x5c7c3315d970, L_0x5c7c3315d970, C4<1>, C4<1>;
v0x5c7c330cabe0_0 .net "in_a", 0 0, L_0x5c7c3315d970;  alias, 1 drivers
v0x5c7c330caca0_0 .net "in_b", 0 0, L_0x5c7c3315d970;  alias, 1 drivers
v0x5c7c330cadf0_0 .net "out", 0 0, L_0x5c7c3315da20;  alias, 1 drivers
S_0x5c7c330cb070 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330c5ee0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330cb810_0 .net "in_a", 0 0, L_0x5c7c3315dc90;  alias, 1 drivers
v0x5c7c330cb8b0_0 .net "out", 0 0, L_0x5c7c3315dd40;  alias, 1 drivers
S_0x5c7c330cb290 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330cb070;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315dd40 .functor NAND 1, L_0x5c7c3315dc90, L_0x5c7c3315dc90, C4<1>, C4<1>;
v0x5c7c330cb500_0 .net "in_a", 0 0, L_0x5c7c3315dc90;  alias, 1 drivers
v0x5c7c330cb5c0_0 .net "in_b", 0 0, L_0x5c7c3315dc90;  alias, 1 drivers
v0x5c7c330cb710_0 .net "out", 0 0, L_0x5c7c3315dd40;  alias, 1 drivers
S_0x5c7c330cc850 .scope module, "mux_gate3" "Mux" 15 10, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330d5bb0_0 .net "in_a", 0 0, L_0x5c7c3315ed50;  1 drivers
v0x5c7c330d5c50_0 .net "in_b", 0 0, L_0x5c7c3315edf0;  1 drivers
v0x5c7c330d5d60_0 .net "out", 0 0, L_0x5c7c3315eb90;  1 drivers
v0x5c7c330d5e00_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330d5ea0_0 .net "sel_out", 0 0, L_0x5c7c3315e080;  1 drivers
v0x5c7c330d6020_0 .net "temp_a_out", 0 0, L_0x5c7c3315e1e0;  1 drivers
v0x5c7c330d61d0_0 .net "temp_b_out", 0 0, L_0x5c7c3315e340;  1 drivers
S_0x5c7c330cca50 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330cc850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330cdab0_0 .net "in_a", 0 0, L_0x5c7c3315ed50;  alias, 1 drivers
v0x5c7c330cdb80_0 .net "in_b", 0 0, L_0x5c7c3315e080;  alias, 1 drivers
v0x5c7c330cdc50_0 .net "out", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
v0x5c7c330cdd70_0 .net "temp_out", 0 0, L_0x5c7c3315e130;  1 drivers
S_0x5c7c330cccc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330cca50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e130 .functor NAND 1, L_0x5c7c3315ed50, L_0x5c7c3315e080, C4<1>, C4<1>;
v0x5c7c330ccf30_0 .net "in_a", 0 0, L_0x5c7c3315ed50;  alias, 1 drivers
v0x5c7c330cd010_0 .net "in_b", 0 0, L_0x5c7c3315e080;  alias, 1 drivers
v0x5c7c330cd0d0_0 .net "out", 0 0, L_0x5c7c3315e130;  alias, 1 drivers
S_0x5c7c330cd1f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330cca50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330cd930_0 .net "in_a", 0 0, L_0x5c7c3315e130;  alias, 1 drivers
v0x5c7c330cd9d0_0 .net "out", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
S_0x5c7c330cd410 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330cd1f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e1e0 .functor NAND 1, L_0x5c7c3315e130, L_0x5c7c3315e130, C4<1>, C4<1>;
v0x5c7c330cd680_0 .net "in_a", 0 0, L_0x5c7c3315e130;  alias, 1 drivers
v0x5c7c330cd740_0 .net "in_b", 0 0, L_0x5c7c3315e130;  alias, 1 drivers
v0x5c7c330cd830_0 .net "out", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
S_0x5c7c330cde30 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330cc850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330cee40_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ceee0_0 .net "in_b", 0 0, L_0x5c7c3315edf0;  alias, 1 drivers
v0x5c7c330cefd0_0 .net "out", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
v0x5c7c330cf0f0_0 .net "temp_out", 0 0, L_0x5c7c3315e290;  1 drivers
S_0x5c7c330ce010 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330cde30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e290 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c3315edf0, C4<1>, C4<1>;
v0x5c7c330ce280_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ce340_0 .net "in_b", 0 0, L_0x5c7c3315edf0;  alias, 1 drivers
v0x5c7c330ce400_0 .net "out", 0 0, L_0x5c7c3315e290;  alias, 1 drivers
S_0x5c7c330ce520 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330cde30;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330cec90_0 .net "in_a", 0 0, L_0x5c7c3315e290;  alias, 1 drivers
v0x5c7c330ced30_0 .net "out", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
S_0x5c7c330ce740 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ce520;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e340 .functor NAND 1, L_0x5c7c3315e290, L_0x5c7c3315e290, C4<1>, C4<1>;
v0x5c7c330ce9b0_0 .net "in_a", 0 0, L_0x5c7c3315e290;  alias, 1 drivers
v0x5c7c330ceaa0_0 .net "in_b", 0 0, L_0x5c7c3315e290;  alias, 1 drivers
v0x5c7c330ceb90_0 .net "out", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
S_0x5c7c330cf1b0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330cc850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330cf8b0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330cf950_0 .net "out", 0 0, L_0x5c7c3315e080;  alias, 1 drivers
S_0x5c7c330cf380 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330cf1b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e080 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330cf5d0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330cf690_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330cf750_0 .net "out", 0 0, L_0x5c7c3315e080;  alias, 1 drivers
S_0x5c7c330cfa50 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330cc850;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330d5500_0 .net "branch1_out", 0 0, L_0x5c7c3315e550;  1 drivers
v0x5c7c330d5630_0 .net "branch2_out", 0 0, L_0x5c7c3315e870;  1 drivers
v0x5c7c330d5780_0 .net "in_a", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
v0x5c7c330d5850_0 .net "in_b", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
v0x5c7c330d58f0_0 .net "out", 0 0, L_0x5c7c3315eb90;  alias, 1 drivers
v0x5c7c330d5990_0 .net "temp1_out", 0 0, L_0x5c7c3315e4a0;  1 drivers
v0x5c7c330d5a30_0 .net "temp2_out", 0 0, L_0x5c7c3315e7c0;  1 drivers
v0x5c7c330d5ad0_0 .net "temp3_out", 0 0, L_0x5c7c3315eae0;  1 drivers
S_0x5c7c330cfc80 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330cfa50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330d0d40_0 .net "in_a", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
v0x5c7c330d0de0_0 .net "in_b", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
v0x5c7c330d0ea0_0 .net "out", 0 0, L_0x5c7c3315e4a0;  alias, 1 drivers
v0x5c7c330d0fc0_0 .net "temp_out", 0 0, L_0x5c7c3315e3f0;  1 drivers
S_0x5c7c330cfef0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330cfc80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e3f0 .functor NAND 1, L_0x5c7c3315e1e0, L_0x5c7c3315e1e0, C4<1>, C4<1>;
v0x5c7c330d0160_0 .net "in_a", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
v0x5c7c330d0220_0 .net "in_b", 0 0, L_0x5c7c3315e1e0;  alias, 1 drivers
v0x5c7c330d0370_0 .net "out", 0 0, L_0x5c7c3315e3f0;  alias, 1 drivers
S_0x5c7c330d0470 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330cfc80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d0b90_0 .net "in_a", 0 0, L_0x5c7c3315e3f0;  alias, 1 drivers
v0x5c7c330d0c30_0 .net "out", 0 0, L_0x5c7c3315e4a0;  alias, 1 drivers
S_0x5c7c330d0640 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d0470;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e4a0 .functor NAND 1, L_0x5c7c3315e3f0, L_0x5c7c3315e3f0, C4<1>, C4<1>;
v0x5c7c330d08b0_0 .net "in_a", 0 0, L_0x5c7c3315e3f0;  alias, 1 drivers
v0x5c7c330d09a0_0 .net "in_b", 0 0, L_0x5c7c3315e3f0;  alias, 1 drivers
v0x5c7c330d0a90_0 .net "out", 0 0, L_0x5c7c3315e4a0;  alias, 1 drivers
S_0x5c7c330d1130 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330cfa50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330d2160_0 .net "in_a", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
v0x5c7c330d2200_0 .net "in_b", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
v0x5c7c330d22c0_0 .net "out", 0 0, L_0x5c7c3315e7c0;  alias, 1 drivers
v0x5c7c330d23e0_0 .net "temp_out", 0 0, L_0x5c7c3315e710;  1 drivers
S_0x5c7c330d1310 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330d1130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e710 .functor NAND 1, L_0x5c7c3315e340, L_0x5c7c3315e340, C4<1>, C4<1>;
v0x5c7c330d1580_0 .net "in_a", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
v0x5c7c330d1640_0 .net "in_b", 0 0, L_0x5c7c3315e340;  alias, 1 drivers
v0x5c7c330d1790_0 .net "out", 0 0, L_0x5c7c3315e710;  alias, 1 drivers
S_0x5c7c330d1890 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330d1130;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d1fb0_0 .net "in_a", 0 0, L_0x5c7c3315e710;  alias, 1 drivers
v0x5c7c330d2050_0 .net "out", 0 0, L_0x5c7c3315e7c0;  alias, 1 drivers
S_0x5c7c330d1a60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d1890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e7c0 .functor NAND 1, L_0x5c7c3315e710, L_0x5c7c3315e710, C4<1>, C4<1>;
v0x5c7c330d1cd0_0 .net "in_a", 0 0, L_0x5c7c3315e710;  alias, 1 drivers
v0x5c7c330d1dc0_0 .net "in_b", 0 0, L_0x5c7c3315e710;  alias, 1 drivers
v0x5c7c330d1eb0_0 .net "out", 0 0, L_0x5c7c3315e7c0;  alias, 1 drivers
S_0x5c7c330d2550 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330cfa50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330d3590_0 .net "in_a", 0 0, L_0x5c7c3315e550;  alias, 1 drivers
v0x5c7c330d3660_0 .net "in_b", 0 0, L_0x5c7c3315e870;  alias, 1 drivers
v0x5c7c330d3730_0 .net "out", 0 0, L_0x5c7c3315eae0;  alias, 1 drivers
v0x5c7c330d3850_0 .net "temp_out", 0 0, L_0x5c7c3315ea30;  1 drivers
S_0x5c7c330d2730 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330d2550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ea30 .functor NAND 1, L_0x5c7c3315e550, L_0x5c7c3315e870, C4<1>, C4<1>;
v0x5c7c330d2980_0 .net "in_a", 0 0, L_0x5c7c3315e550;  alias, 1 drivers
v0x5c7c330d2a60_0 .net "in_b", 0 0, L_0x5c7c3315e870;  alias, 1 drivers
v0x5c7c330d2b20_0 .net "out", 0 0, L_0x5c7c3315ea30;  alias, 1 drivers
S_0x5c7c330d2c70 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330d2550;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d33e0_0 .net "in_a", 0 0, L_0x5c7c3315ea30;  alias, 1 drivers
v0x5c7c330d3480_0 .net "out", 0 0, L_0x5c7c3315eae0;  alias, 1 drivers
S_0x5c7c330d2e90 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d2c70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315eae0 .functor NAND 1, L_0x5c7c3315ea30, L_0x5c7c3315ea30, C4<1>, C4<1>;
v0x5c7c330d3100_0 .net "in_a", 0 0, L_0x5c7c3315ea30;  alias, 1 drivers
v0x5c7c330d31f0_0 .net "in_b", 0 0, L_0x5c7c3315ea30;  alias, 1 drivers
v0x5c7c330d32e0_0 .net "out", 0 0, L_0x5c7c3315eae0;  alias, 1 drivers
S_0x5c7c330d39a0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330cfa50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d40d0_0 .net "in_a", 0 0, L_0x5c7c3315e4a0;  alias, 1 drivers
v0x5c7c330d4170_0 .net "out", 0 0, L_0x5c7c3315e550;  alias, 1 drivers
S_0x5c7c330d3b70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d39a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e550 .functor NAND 1, L_0x5c7c3315e4a0, L_0x5c7c3315e4a0, C4<1>, C4<1>;
v0x5c7c330d3de0_0 .net "in_a", 0 0, L_0x5c7c3315e4a0;  alias, 1 drivers
v0x5c7c330d3ea0_0 .net "in_b", 0 0, L_0x5c7c3315e4a0;  alias, 1 drivers
v0x5c7c330d3ff0_0 .net "out", 0 0, L_0x5c7c3315e550;  alias, 1 drivers
S_0x5c7c330d4270 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330cfa50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d4a40_0 .net "in_a", 0 0, L_0x5c7c3315e7c0;  alias, 1 drivers
v0x5c7c330d4ae0_0 .net "out", 0 0, L_0x5c7c3315e870;  alias, 1 drivers
S_0x5c7c330d44e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d4270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315e870 .functor NAND 1, L_0x5c7c3315e7c0, L_0x5c7c3315e7c0, C4<1>, C4<1>;
v0x5c7c330d4750_0 .net "in_a", 0 0, L_0x5c7c3315e7c0;  alias, 1 drivers
v0x5c7c330d4810_0 .net "in_b", 0 0, L_0x5c7c3315e7c0;  alias, 1 drivers
v0x5c7c330d4960_0 .net "out", 0 0, L_0x5c7c3315e870;  alias, 1 drivers
S_0x5c7c330d4be0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330cfa50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d5380_0 .net "in_a", 0 0, L_0x5c7c3315eae0;  alias, 1 drivers
v0x5c7c330d5420_0 .net "out", 0 0, L_0x5c7c3315eb90;  alias, 1 drivers
S_0x5c7c330d4e00 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d4be0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315eb90 .functor NAND 1, L_0x5c7c3315eae0, L_0x5c7c3315eae0, C4<1>, C4<1>;
v0x5c7c330d5070_0 .net "in_a", 0 0, L_0x5c7c3315eae0;  alias, 1 drivers
v0x5c7c330d5130_0 .net "in_b", 0 0, L_0x5c7c3315eae0;  alias, 1 drivers
v0x5c7c330d5280_0 .net "out", 0 0, L_0x5c7c3315eb90;  alias, 1 drivers
S_0x5c7c330d63c0 .scope module, "mux_gate4" "Mux" 15 11, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330dff30_0 .net "in_a", 0 0, L_0x5c7c3315fb60;  1 drivers
v0x5c7c330dffd0_0 .net "in_b", 0 0, L_0x5c7c3315fd10;  1 drivers
v0x5c7c330e00e0_0 .net "out", 0 0, L_0x5c7c3315f9a0;  1 drivers
v0x5c7c330e0180_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e0220_0 .net "sel_out", 0 0, L_0x5c7c3315ee90;  1 drivers
v0x5c7c330e03a0_0 .net "temp_a_out", 0 0, L_0x5c7c3315eff0;  1 drivers
v0x5c7c330e0550_0 .net "temp_b_out", 0 0, L_0x5c7c3315f150;  1 drivers
S_0x5c7c330d65c0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330d63c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330d7620_0 .net "in_a", 0 0, L_0x5c7c3315fb60;  alias, 1 drivers
v0x5c7c330d76f0_0 .net "in_b", 0 0, L_0x5c7c3315ee90;  alias, 1 drivers
v0x5c7c330d77c0_0 .net "out", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
v0x5c7c330d78e0_0 .net "temp_out", 0 0, L_0x5c7c3315ef40;  1 drivers
S_0x5c7c330d6830 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330d65c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ef40 .functor NAND 1, L_0x5c7c3315fb60, L_0x5c7c3315ee90, C4<1>, C4<1>;
v0x5c7c330d6aa0_0 .net "in_a", 0 0, L_0x5c7c3315fb60;  alias, 1 drivers
v0x5c7c330d6b80_0 .net "in_b", 0 0, L_0x5c7c3315ee90;  alias, 1 drivers
v0x5c7c330d6c40_0 .net "out", 0 0, L_0x5c7c3315ef40;  alias, 1 drivers
S_0x5c7c330d6d60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330d65c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d74a0_0 .net "in_a", 0 0, L_0x5c7c3315ef40;  alias, 1 drivers
v0x5c7c330d7540_0 .net "out", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
S_0x5c7c330d6f80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d6d60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315eff0 .functor NAND 1, L_0x5c7c3315ef40, L_0x5c7c3315ef40, C4<1>, C4<1>;
v0x5c7c330d71f0_0 .net "in_a", 0 0, L_0x5c7c3315ef40;  alias, 1 drivers
v0x5c7c330d72b0_0 .net "in_b", 0 0, L_0x5c7c3315ef40;  alias, 1 drivers
v0x5c7c330d73a0_0 .net "out", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
S_0x5c7c330d79a0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330d63c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330d89b0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330d8a50_0 .net "in_b", 0 0, L_0x5c7c3315fd10;  alias, 1 drivers
v0x5c7c330d8b40_0 .net "out", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
v0x5c7c330d8c60_0 .net "temp_out", 0 0, L_0x5c7c3315f0a0;  1 drivers
S_0x5c7c330d7b80 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330d79a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f0a0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c3315fd10, C4<1>, C4<1>;
v0x5c7c330d7df0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330d7eb0_0 .net "in_b", 0 0, L_0x5c7c3315fd10;  alias, 1 drivers
v0x5c7c330d7f70_0 .net "out", 0 0, L_0x5c7c3315f0a0;  alias, 1 drivers
S_0x5c7c330d8090 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330d79a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d8800_0 .net "in_a", 0 0, L_0x5c7c3315f0a0;  alias, 1 drivers
v0x5c7c330d88a0_0 .net "out", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
S_0x5c7c330d82b0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d8090;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f150 .functor NAND 1, L_0x5c7c3315f0a0, L_0x5c7c3315f0a0, C4<1>, C4<1>;
v0x5c7c330d8520_0 .net "in_a", 0 0, L_0x5c7c3315f0a0;  alias, 1 drivers
v0x5c7c330d8610_0 .net "in_b", 0 0, L_0x5c7c3315f0a0;  alias, 1 drivers
v0x5c7c330d8700_0 .net "out", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
S_0x5c7c330d8d20 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330d63c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330d9420_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330d9cd0_0 .net "out", 0 0, L_0x5c7c3315ee90;  alias, 1 drivers
S_0x5c7c330d8ef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330d8d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ee90 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330d9140_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330d9200_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330d92c0_0 .net "out", 0 0, L_0x5c7c3315ee90;  alias, 1 drivers
S_0x5c7c330d9dd0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330d63c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330df880_0 .net "branch1_out", 0 0, L_0x5c7c3315f360;  1 drivers
v0x5c7c330df9b0_0 .net "branch2_out", 0 0, L_0x5c7c3315f680;  1 drivers
v0x5c7c330dfb00_0 .net "in_a", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
v0x5c7c330dfbd0_0 .net "in_b", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
v0x5c7c330dfc70_0 .net "out", 0 0, L_0x5c7c3315f9a0;  alias, 1 drivers
v0x5c7c330dfd10_0 .net "temp1_out", 0 0, L_0x5c7c3315f2b0;  1 drivers
v0x5c7c330dfdb0_0 .net "temp2_out", 0 0, L_0x5c7c3315f5d0;  1 drivers
v0x5c7c330dfe50_0 .net "temp3_out", 0 0, L_0x5c7c3315f8f0;  1 drivers
S_0x5c7c330da000 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330d9dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330db0c0_0 .net "in_a", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
v0x5c7c330db160_0 .net "in_b", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
v0x5c7c330db220_0 .net "out", 0 0, L_0x5c7c3315f2b0;  alias, 1 drivers
v0x5c7c330db340_0 .net "temp_out", 0 0, L_0x5c7c3315f200;  1 drivers
S_0x5c7c330da270 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330da000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f200 .functor NAND 1, L_0x5c7c3315eff0, L_0x5c7c3315eff0, C4<1>, C4<1>;
v0x5c7c330da4e0_0 .net "in_a", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
v0x5c7c330da5a0_0 .net "in_b", 0 0, L_0x5c7c3315eff0;  alias, 1 drivers
v0x5c7c330da6f0_0 .net "out", 0 0, L_0x5c7c3315f200;  alias, 1 drivers
S_0x5c7c330da7f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330da000;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330daf10_0 .net "in_a", 0 0, L_0x5c7c3315f200;  alias, 1 drivers
v0x5c7c330dafb0_0 .net "out", 0 0, L_0x5c7c3315f2b0;  alias, 1 drivers
S_0x5c7c330da9c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330da7f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f2b0 .functor NAND 1, L_0x5c7c3315f200, L_0x5c7c3315f200, C4<1>, C4<1>;
v0x5c7c330dac30_0 .net "in_a", 0 0, L_0x5c7c3315f200;  alias, 1 drivers
v0x5c7c330dad20_0 .net "in_b", 0 0, L_0x5c7c3315f200;  alias, 1 drivers
v0x5c7c330dae10_0 .net "out", 0 0, L_0x5c7c3315f2b0;  alias, 1 drivers
S_0x5c7c330db4b0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330d9dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330dc4e0_0 .net "in_a", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
v0x5c7c330dc580_0 .net "in_b", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
v0x5c7c330dc640_0 .net "out", 0 0, L_0x5c7c3315f5d0;  alias, 1 drivers
v0x5c7c330dc760_0 .net "temp_out", 0 0, L_0x5c7c3315f520;  1 drivers
S_0x5c7c330db690 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330db4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f520 .functor NAND 1, L_0x5c7c3315f150, L_0x5c7c3315f150, C4<1>, C4<1>;
v0x5c7c330db900_0 .net "in_a", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
v0x5c7c330db9c0_0 .net "in_b", 0 0, L_0x5c7c3315f150;  alias, 1 drivers
v0x5c7c330dbb10_0 .net "out", 0 0, L_0x5c7c3315f520;  alias, 1 drivers
S_0x5c7c330dbc10 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330db4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330dc330_0 .net "in_a", 0 0, L_0x5c7c3315f520;  alias, 1 drivers
v0x5c7c330dc3d0_0 .net "out", 0 0, L_0x5c7c3315f5d0;  alias, 1 drivers
S_0x5c7c330dbde0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330dbc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f5d0 .functor NAND 1, L_0x5c7c3315f520, L_0x5c7c3315f520, C4<1>, C4<1>;
v0x5c7c330dc050_0 .net "in_a", 0 0, L_0x5c7c3315f520;  alias, 1 drivers
v0x5c7c330dc140_0 .net "in_b", 0 0, L_0x5c7c3315f520;  alias, 1 drivers
v0x5c7c330dc230_0 .net "out", 0 0, L_0x5c7c3315f5d0;  alias, 1 drivers
S_0x5c7c330dc8d0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330d9dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330dd910_0 .net "in_a", 0 0, L_0x5c7c3315f360;  alias, 1 drivers
v0x5c7c330dd9e0_0 .net "in_b", 0 0, L_0x5c7c3315f680;  alias, 1 drivers
v0x5c7c330ddab0_0 .net "out", 0 0, L_0x5c7c3315f8f0;  alias, 1 drivers
v0x5c7c330ddbd0_0 .net "temp_out", 0 0, L_0x5c7c3315f840;  1 drivers
S_0x5c7c330dcab0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330dc8d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f840 .functor NAND 1, L_0x5c7c3315f360, L_0x5c7c3315f680, C4<1>, C4<1>;
v0x5c7c330dcd00_0 .net "in_a", 0 0, L_0x5c7c3315f360;  alias, 1 drivers
v0x5c7c330dcde0_0 .net "in_b", 0 0, L_0x5c7c3315f680;  alias, 1 drivers
v0x5c7c330dcea0_0 .net "out", 0 0, L_0x5c7c3315f840;  alias, 1 drivers
S_0x5c7c330dcff0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330dc8d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330dd760_0 .net "in_a", 0 0, L_0x5c7c3315f840;  alias, 1 drivers
v0x5c7c330dd800_0 .net "out", 0 0, L_0x5c7c3315f8f0;  alias, 1 drivers
S_0x5c7c330dd210 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330dcff0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f8f0 .functor NAND 1, L_0x5c7c3315f840, L_0x5c7c3315f840, C4<1>, C4<1>;
v0x5c7c330dd480_0 .net "in_a", 0 0, L_0x5c7c3315f840;  alias, 1 drivers
v0x5c7c330dd570_0 .net "in_b", 0 0, L_0x5c7c3315f840;  alias, 1 drivers
v0x5c7c330dd660_0 .net "out", 0 0, L_0x5c7c3315f8f0;  alias, 1 drivers
S_0x5c7c330ddd20 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330d9dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330de450_0 .net "in_a", 0 0, L_0x5c7c3315f2b0;  alias, 1 drivers
v0x5c7c330de4f0_0 .net "out", 0 0, L_0x5c7c3315f360;  alias, 1 drivers
S_0x5c7c330ddef0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ddd20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f360 .functor NAND 1, L_0x5c7c3315f2b0, L_0x5c7c3315f2b0, C4<1>, C4<1>;
v0x5c7c330de160_0 .net "in_a", 0 0, L_0x5c7c3315f2b0;  alias, 1 drivers
v0x5c7c330de220_0 .net "in_b", 0 0, L_0x5c7c3315f2b0;  alias, 1 drivers
v0x5c7c330de370_0 .net "out", 0 0, L_0x5c7c3315f360;  alias, 1 drivers
S_0x5c7c330de5f0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330d9dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330dedc0_0 .net "in_a", 0 0, L_0x5c7c3315f5d0;  alias, 1 drivers
v0x5c7c330dee60_0 .net "out", 0 0, L_0x5c7c3315f680;  alias, 1 drivers
S_0x5c7c330de860 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330de5f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f680 .functor NAND 1, L_0x5c7c3315f5d0, L_0x5c7c3315f5d0, C4<1>, C4<1>;
v0x5c7c330dead0_0 .net "in_a", 0 0, L_0x5c7c3315f5d0;  alias, 1 drivers
v0x5c7c330deb90_0 .net "in_b", 0 0, L_0x5c7c3315f5d0;  alias, 1 drivers
v0x5c7c330dece0_0 .net "out", 0 0, L_0x5c7c3315f680;  alias, 1 drivers
S_0x5c7c330def60 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330d9dd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330df700_0 .net "in_a", 0 0, L_0x5c7c3315f8f0;  alias, 1 drivers
v0x5c7c330df7a0_0 .net "out", 0 0, L_0x5c7c3315f9a0;  alias, 1 drivers
S_0x5c7c330df180 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330def60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315f9a0 .functor NAND 1, L_0x5c7c3315f8f0, L_0x5c7c3315f8f0, C4<1>, C4<1>;
v0x5c7c330df3f0_0 .net "in_a", 0 0, L_0x5c7c3315f8f0;  alias, 1 drivers
v0x5c7c330df4b0_0 .net "in_b", 0 0, L_0x5c7c3315f8f0;  alias, 1 drivers
v0x5c7c330df600_0 .net "out", 0 0, L_0x5c7c3315f9a0;  alias, 1 drivers
S_0x5c7c330e0740 .scope module, "mux_gate5" "Mux" 15 12, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330e9aa0_0 .net "in_a", 0 0, L_0x5c7c33160bf0;  1 drivers
v0x5c7c330e9b40_0 .net "in_b", 0 0, L_0x5c7c33160c90;  1 drivers
v0x5c7c330e9c50_0 .net "out", 0 0, L_0x5c7c33160a30;  1 drivers
v0x5c7c330e9cf0_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e9d90_0 .net "sel_out", 0 0, L_0x5c7c3315ff20;  1 drivers
v0x5c7c330e9f10_0 .net "temp_a_out", 0 0, L_0x5c7c33160080;  1 drivers
v0x5c7c330ea0c0_0 .net "temp_b_out", 0 0, L_0x5c7c331601e0;  1 drivers
S_0x5c7c330e0940 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330e0740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330e19a0_0 .net "in_a", 0 0, L_0x5c7c33160bf0;  alias, 1 drivers
v0x5c7c330e1a70_0 .net "in_b", 0 0, L_0x5c7c3315ff20;  alias, 1 drivers
v0x5c7c330e1b40_0 .net "out", 0 0, L_0x5c7c33160080;  alias, 1 drivers
v0x5c7c330e1c60_0 .net "temp_out", 0 0, L_0x5c7c3315ffd0;  1 drivers
S_0x5c7c330e0bb0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330e0940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ffd0 .functor NAND 1, L_0x5c7c33160bf0, L_0x5c7c3315ff20, C4<1>, C4<1>;
v0x5c7c330e0e20_0 .net "in_a", 0 0, L_0x5c7c33160bf0;  alias, 1 drivers
v0x5c7c330e0f00_0 .net "in_b", 0 0, L_0x5c7c3315ff20;  alias, 1 drivers
v0x5c7c330e0fc0_0 .net "out", 0 0, L_0x5c7c3315ffd0;  alias, 1 drivers
S_0x5c7c330e10e0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330e0940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e1820_0 .net "in_a", 0 0, L_0x5c7c3315ffd0;  alias, 1 drivers
v0x5c7c330e18c0_0 .net "out", 0 0, L_0x5c7c33160080;  alias, 1 drivers
S_0x5c7c330e1300 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e10e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160080 .functor NAND 1, L_0x5c7c3315ffd0, L_0x5c7c3315ffd0, C4<1>, C4<1>;
v0x5c7c330e1570_0 .net "in_a", 0 0, L_0x5c7c3315ffd0;  alias, 1 drivers
v0x5c7c330e1630_0 .net "in_b", 0 0, L_0x5c7c3315ffd0;  alias, 1 drivers
v0x5c7c330e1720_0 .net "out", 0 0, L_0x5c7c33160080;  alias, 1 drivers
S_0x5c7c330e1d20 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330e0740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330e2d30_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e2dd0_0 .net "in_b", 0 0, L_0x5c7c33160c90;  alias, 1 drivers
v0x5c7c330e2ec0_0 .net "out", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
v0x5c7c330e2fe0_0 .net "temp_out", 0 0, L_0x5c7c33160130;  1 drivers
S_0x5c7c330e1f00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330e1d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160130 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33160c90, C4<1>, C4<1>;
v0x5c7c330e2170_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e2230_0 .net "in_b", 0 0, L_0x5c7c33160c90;  alias, 1 drivers
v0x5c7c330e22f0_0 .net "out", 0 0, L_0x5c7c33160130;  alias, 1 drivers
S_0x5c7c330e2410 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330e1d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e2b80_0 .net "in_a", 0 0, L_0x5c7c33160130;  alias, 1 drivers
v0x5c7c330e2c20_0 .net "out", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
S_0x5c7c330e2630 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e2410;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331601e0 .functor NAND 1, L_0x5c7c33160130, L_0x5c7c33160130, C4<1>, C4<1>;
v0x5c7c330e28a0_0 .net "in_a", 0 0, L_0x5c7c33160130;  alias, 1 drivers
v0x5c7c330e2990_0 .net "in_b", 0 0, L_0x5c7c33160130;  alias, 1 drivers
v0x5c7c330e2a80_0 .net "out", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
S_0x5c7c330e30a0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330e0740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e37a0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e3840_0 .net "out", 0 0, L_0x5c7c3315ff20;  alias, 1 drivers
S_0x5c7c330e3270 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e30a0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c3315ff20 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330e34c0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e3580_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330e3640_0 .net "out", 0 0, L_0x5c7c3315ff20;  alias, 1 drivers
S_0x5c7c330e3940 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330e0740;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330e93f0_0 .net "branch1_out", 0 0, L_0x5c7c331603f0;  1 drivers
v0x5c7c330e9520_0 .net "branch2_out", 0 0, L_0x5c7c33160710;  1 drivers
v0x5c7c330e9670_0 .net "in_a", 0 0, L_0x5c7c33160080;  alias, 1 drivers
v0x5c7c330e9740_0 .net "in_b", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
v0x5c7c330e97e0_0 .net "out", 0 0, L_0x5c7c33160a30;  alias, 1 drivers
v0x5c7c330e9880_0 .net "temp1_out", 0 0, L_0x5c7c33160340;  1 drivers
v0x5c7c330e9920_0 .net "temp2_out", 0 0, L_0x5c7c33160660;  1 drivers
v0x5c7c330e99c0_0 .net "temp3_out", 0 0, L_0x5c7c33160980;  1 drivers
S_0x5c7c330e3b70 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330e3940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330e4c30_0 .net "in_a", 0 0, L_0x5c7c33160080;  alias, 1 drivers
v0x5c7c330e4cd0_0 .net "in_b", 0 0, L_0x5c7c33160080;  alias, 1 drivers
v0x5c7c330e4d90_0 .net "out", 0 0, L_0x5c7c33160340;  alias, 1 drivers
v0x5c7c330e4eb0_0 .net "temp_out", 0 0, L_0x5c7c33160290;  1 drivers
S_0x5c7c330e3de0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330e3b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160290 .functor NAND 1, L_0x5c7c33160080, L_0x5c7c33160080, C4<1>, C4<1>;
v0x5c7c330e4050_0 .net "in_a", 0 0, L_0x5c7c33160080;  alias, 1 drivers
v0x5c7c330e4110_0 .net "in_b", 0 0, L_0x5c7c33160080;  alias, 1 drivers
v0x5c7c330e4260_0 .net "out", 0 0, L_0x5c7c33160290;  alias, 1 drivers
S_0x5c7c330e4360 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330e3b70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e4a80_0 .net "in_a", 0 0, L_0x5c7c33160290;  alias, 1 drivers
v0x5c7c330e4b20_0 .net "out", 0 0, L_0x5c7c33160340;  alias, 1 drivers
S_0x5c7c330e4530 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e4360;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160340 .functor NAND 1, L_0x5c7c33160290, L_0x5c7c33160290, C4<1>, C4<1>;
v0x5c7c330e47a0_0 .net "in_a", 0 0, L_0x5c7c33160290;  alias, 1 drivers
v0x5c7c330e4890_0 .net "in_b", 0 0, L_0x5c7c33160290;  alias, 1 drivers
v0x5c7c330e4980_0 .net "out", 0 0, L_0x5c7c33160340;  alias, 1 drivers
S_0x5c7c330e5020 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330e3940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330e6050_0 .net "in_a", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
v0x5c7c330e60f0_0 .net "in_b", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
v0x5c7c330e61b0_0 .net "out", 0 0, L_0x5c7c33160660;  alias, 1 drivers
v0x5c7c330e62d0_0 .net "temp_out", 0 0, L_0x5c7c331605b0;  1 drivers
S_0x5c7c330e5200 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330e5020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331605b0 .functor NAND 1, L_0x5c7c331601e0, L_0x5c7c331601e0, C4<1>, C4<1>;
v0x5c7c330e5470_0 .net "in_a", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
v0x5c7c330e5530_0 .net "in_b", 0 0, L_0x5c7c331601e0;  alias, 1 drivers
v0x5c7c330e5680_0 .net "out", 0 0, L_0x5c7c331605b0;  alias, 1 drivers
S_0x5c7c330e5780 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330e5020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e5ea0_0 .net "in_a", 0 0, L_0x5c7c331605b0;  alias, 1 drivers
v0x5c7c330e5f40_0 .net "out", 0 0, L_0x5c7c33160660;  alias, 1 drivers
S_0x5c7c330e5950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e5780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160660 .functor NAND 1, L_0x5c7c331605b0, L_0x5c7c331605b0, C4<1>, C4<1>;
v0x5c7c330e5bc0_0 .net "in_a", 0 0, L_0x5c7c331605b0;  alias, 1 drivers
v0x5c7c330e5cb0_0 .net "in_b", 0 0, L_0x5c7c331605b0;  alias, 1 drivers
v0x5c7c330e5da0_0 .net "out", 0 0, L_0x5c7c33160660;  alias, 1 drivers
S_0x5c7c330e6440 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330e3940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330e7480_0 .net "in_a", 0 0, L_0x5c7c331603f0;  alias, 1 drivers
v0x5c7c330e7550_0 .net "in_b", 0 0, L_0x5c7c33160710;  alias, 1 drivers
v0x5c7c330e7620_0 .net "out", 0 0, L_0x5c7c33160980;  alias, 1 drivers
v0x5c7c330e7740_0 .net "temp_out", 0 0, L_0x5c7c331608d0;  1 drivers
S_0x5c7c330e6620 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330e6440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331608d0 .functor NAND 1, L_0x5c7c331603f0, L_0x5c7c33160710, C4<1>, C4<1>;
v0x5c7c330e6870_0 .net "in_a", 0 0, L_0x5c7c331603f0;  alias, 1 drivers
v0x5c7c330e6950_0 .net "in_b", 0 0, L_0x5c7c33160710;  alias, 1 drivers
v0x5c7c330e6a10_0 .net "out", 0 0, L_0x5c7c331608d0;  alias, 1 drivers
S_0x5c7c330e6b60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330e6440;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e72d0_0 .net "in_a", 0 0, L_0x5c7c331608d0;  alias, 1 drivers
v0x5c7c330e7370_0 .net "out", 0 0, L_0x5c7c33160980;  alias, 1 drivers
S_0x5c7c330e6d80 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e6b60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160980 .functor NAND 1, L_0x5c7c331608d0, L_0x5c7c331608d0, C4<1>, C4<1>;
v0x5c7c330e6ff0_0 .net "in_a", 0 0, L_0x5c7c331608d0;  alias, 1 drivers
v0x5c7c330e70e0_0 .net "in_b", 0 0, L_0x5c7c331608d0;  alias, 1 drivers
v0x5c7c330e71d0_0 .net "out", 0 0, L_0x5c7c33160980;  alias, 1 drivers
S_0x5c7c330e7890 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330e3940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e7fc0_0 .net "in_a", 0 0, L_0x5c7c33160340;  alias, 1 drivers
v0x5c7c330e8060_0 .net "out", 0 0, L_0x5c7c331603f0;  alias, 1 drivers
S_0x5c7c330e7a60 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e7890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331603f0 .functor NAND 1, L_0x5c7c33160340, L_0x5c7c33160340, C4<1>, C4<1>;
v0x5c7c330e7cd0_0 .net "in_a", 0 0, L_0x5c7c33160340;  alias, 1 drivers
v0x5c7c330e7d90_0 .net "in_b", 0 0, L_0x5c7c33160340;  alias, 1 drivers
v0x5c7c330e7ee0_0 .net "out", 0 0, L_0x5c7c331603f0;  alias, 1 drivers
S_0x5c7c330e8160 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330e3940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e8930_0 .net "in_a", 0 0, L_0x5c7c33160660;  alias, 1 drivers
v0x5c7c330e89d0_0 .net "out", 0 0, L_0x5c7c33160710;  alias, 1 drivers
S_0x5c7c330e83d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e8160;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160710 .functor NAND 1, L_0x5c7c33160660, L_0x5c7c33160660, C4<1>, C4<1>;
v0x5c7c330e8640_0 .net "in_a", 0 0, L_0x5c7c33160660;  alias, 1 drivers
v0x5c7c330e8700_0 .net "in_b", 0 0, L_0x5c7c33160660;  alias, 1 drivers
v0x5c7c330e8850_0 .net "out", 0 0, L_0x5c7c33160710;  alias, 1 drivers
S_0x5c7c330e8ad0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330e3940;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330e9270_0 .net "in_a", 0 0, L_0x5c7c33160980;  alias, 1 drivers
v0x5c7c330e9310_0 .net "out", 0 0, L_0x5c7c33160a30;  alias, 1 drivers
S_0x5c7c330e8cf0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330e8ad0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160a30 .functor NAND 1, L_0x5c7c33160980, L_0x5c7c33160980, C4<1>, C4<1>;
v0x5c7c330e8f60_0 .net "in_a", 0 0, L_0x5c7c33160980;  alias, 1 drivers
v0x5c7c330e9020_0 .net "in_b", 0 0, L_0x5c7c33160980;  alias, 1 drivers
v0x5c7c330e9170_0 .net "out", 0 0, L_0x5c7c33160a30;  alias, 1 drivers
S_0x5c7c330ea2b0 .scope module, "mux_gate6" "Mux" 15 13, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330f3610_0 .net "in_a", 0 0, L_0x5c7c33161a70;  1 drivers
v0x5c7c330f36b0_0 .net "in_b", 0 0, L_0x5c7c33161b10;  1 drivers
v0x5c7c330f37c0_0 .net "out", 0 0, L_0x5c7c331618b0;  1 drivers
v0x5c7c330f3860_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330f3900_0 .net "sel_out", 0 0, L_0x5c7c33160da0;  1 drivers
v0x5c7c330f3a80_0 .net "temp_a_out", 0 0, L_0x5c7c33160f00;  1 drivers
v0x5c7c330f3c30_0 .net "temp_b_out", 0 0, L_0x5c7c33161060;  1 drivers
S_0x5c7c330ea4b0 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330ea2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330eb510_0 .net "in_a", 0 0, L_0x5c7c33161a70;  alias, 1 drivers
v0x5c7c330eb5e0_0 .net "in_b", 0 0, L_0x5c7c33160da0;  alias, 1 drivers
v0x5c7c330eb6b0_0 .net "out", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
v0x5c7c330eb7d0_0 .net "temp_out", 0 0, L_0x5c7c33160e50;  1 drivers
S_0x5c7c330ea720 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330ea4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160e50 .functor NAND 1, L_0x5c7c33161a70, L_0x5c7c33160da0, C4<1>, C4<1>;
v0x5c7c330ea990_0 .net "in_a", 0 0, L_0x5c7c33161a70;  alias, 1 drivers
v0x5c7c330eaa70_0 .net "in_b", 0 0, L_0x5c7c33160da0;  alias, 1 drivers
v0x5c7c330eab30_0 .net "out", 0 0, L_0x5c7c33160e50;  alias, 1 drivers
S_0x5c7c330eac50 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330ea4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330eb390_0 .net "in_a", 0 0, L_0x5c7c33160e50;  alias, 1 drivers
v0x5c7c330eb430_0 .net "out", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
S_0x5c7c330eae70 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330eac50;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160f00 .functor NAND 1, L_0x5c7c33160e50, L_0x5c7c33160e50, C4<1>, C4<1>;
v0x5c7c330eb0e0_0 .net "in_a", 0 0, L_0x5c7c33160e50;  alias, 1 drivers
v0x5c7c330eb1a0_0 .net "in_b", 0 0, L_0x5c7c33160e50;  alias, 1 drivers
v0x5c7c330eb290_0 .net "out", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
S_0x5c7c330eb890 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330ea2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330ec8a0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ec940_0 .net "in_b", 0 0, L_0x5c7c33161b10;  alias, 1 drivers
v0x5c7c330eca30_0 .net "out", 0 0, L_0x5c7c33161060;  alias, 1 drivers
v0x5c7c330ecb50_0 .net "temp_out", 0 0, L_0x5c7c33160fb0;  1 drivers
S_0x5c7c330eba70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330eb890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160fb0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33161b10, C4<1>, C4<1>;
v0x5c7c330ebce0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ebda0_0 .net "in_b", 0 0, L_0x5c7c33161b10;  alias, 1 drivers
v0x5c7c330ebe60_0 .net "out", 0 0, L_0x5c7c33160fb0;  alias, 1 drivers
S_0x5c7c330ebf80 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330eb890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ec6f0_0 .net "in_a", 0 0, L_0x5c7c33160fb0;  alias, 1 drivers
v0x5c7c330ec790_0 .net "out", 0 0, L_0x5c7c33161060;  alias, 1 drivers
S_0x5c7c330ec1a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ebf80;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161060 .functor NAND 1, L_0x5c7c33160fb0, L_0x5c7c33160fb0, C4<1>, C4<1>;
v0x5c7c330ec410_0 .net "in_a", 0 0, L_0x5c7c33160fb0;  alias, 1 drivers
v0x5c7c330ec500_0 .net "in_b", 0 0, L_0x5c7c33160fb0;  alias, 1 drivers
v0x5c7c330ec5f0_0 .net "out", 0 0, L_0x5c7c33161060;  alias, 1 drivers
S_0x5c7c330ecc10 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330ea2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ed310_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ed3b0_0 .net "out", 0 0, L_0x5c7c33160da0;  alias, 1 drivers
S_0x5c7c330ecde0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ecc10;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160da0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330ed030_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ed0f0_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ed1b0_0 .net "out", 0 0, L_0x5c7c33160da0;  alias, 1 drivers
S_0x5c7c330ed4b0 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330ea2b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330f2f60_0 .net "branch1_out", 0 0, L_0x5c7c33161270;  1 drivers
v0x5c7c330f3090_0 .net "branch2_out", 0 0, L_0x5c7c33161590;  1 drivers
v0x5c7c330f31e0_0 .net "in_a", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
v0x5c7c330f32b0_0 .net "in_b", 0 0, L_0x5c7c33161060;  alias, 1 drivers
v0x5c7c330f3350_0 .net "out", 0 0, L_0x5c7c331618b0;  alias, 1 drivers
v0x5c7c330f33f0_0 .net "temp1_out", 0 0, L_0x5c7c331611c0;  1 drivers
v0x5c7c330f3490_0 .net "temp2_out", 0 0, L_0x5c7c331614e0;  1 drivers
v0x5c7c330f3530_0 .net "temp3_out", 0 0, L_0x5c7c33161800;  1 drivers
S_0x5c7c330ed6e0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330ed4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330ee7a0_0 .net "in_a", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
v0x5c7c330ee840_0 .net "in_b", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
v0x5c7c330ee900_0 .net "out", 0 0, L_0x5c7c331611c0;  alias, 1 drivers
v0x5c7c330eea20_0 .net "temp_out", 0 0, L_0x5c7c33161110;  1 drivers
S_0x5c7c330ed950 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330ed6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161110 .functor NAND 1, L_0x5c7c33160f00, L_0x5c7c33160f00, C4<1>, C4<1>;
v0x5c7c330edbc0_0 .net "in_a", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
v0x5c7c330edc80_0 .net "in_b", 0 0, L_0x5c7c33160f00;  alias, 1 drivers
v0x5c7c330eddd0_0 .net "out", 0 0, L_0x5c7c33161110;  alias, 1 drivers
S_0x5c7c330eded0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330ed6e0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ee5f0_0 .net "in_a", 0 0, L_0x5c7c33161110;  alias, 1 drivers
v0x5c7c330ee690_0 .net "out", 0 0, L_0x5c7c331611c0;  alias, 1 drivers
S_0x5c7c330ee0a0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330eded0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331611c0 .functor NAND 1, L_0x5c7c33161110, L_0x5c7c33161110, C4<1>, C4<1>;
v0x5c7c330ee310_0 .net "in_a", 0 0, L_0x5c7c33161110;  alias, 1 drivers
v0x5c7c330ee400_0 .net "in_b", 0 0, L_0x5c7c33161110;  alias, 1 drivers
v0x5c7c330ee4f0_0 .net "out", 0 0, L_0x5c7c331611c0;  alias, 1 drivers
S_0x5c7c330eeb90 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330ed4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330efbc0_0 .net "in_a", 0 0, L_0x5c7c33161060;  alias, 1 drivers
v0x5c7c330efc60_0 .net "in_b", 0 0, L_0x5c7c33161060;  alias, 1 drivers
v0x5c7c330efd20_0 .net "out", 0 0, L_0x5c7c331614e0;  alias, 1 drivers
v0x5c7c330efe40_0 .net "temp_out", 0 0, L_0x5c7c33161430;  1 drivers
S_0x5c7c330eed70 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330eeb90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161430 .functor NAND 1, L_0x5c7c33161060, L_0x5c7c33161060, C4<1>, C4<1>;
v0x5c7c330eefe0_0 .net "in_a", 0 0, L_0x5c7c33161060;  alias, 1 drivers
v0x5c7c330ef0a0_0 .net "in_b", 0 0, L_0x5c7c33161060;  alias, 1 drivers
v0x5c7c330ef1f0_0 .net "out", 0 0, L_0x5c7c33161430;  alias, 1 drivers
S_0x5c7c330ef2f0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330eeb90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330efa10_0 .net "in_a", 0 0, L_0x5c7c33161430;  alias, 1 drivers
v0x5c7c330efab0_0 .net "out", 0 0, L_0x5c7c331614e0;  alias, 1 drivers
S_0x5c7c330ef4c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ef2f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331614e0 .functor NAND 1, L_0x5c7c33161430, L_0x5c7c33161430, C4<1>, C4<1>;
v0x5c7c330ef730_0 .net "in_a", 0 0, L_0x5c7c33161430;  alias, 1 drivers
v0x5c7c330ef820_0 .net "in_b", 0 0, L_0x5c7c33161430;  alias, 1 drivers
v0x5c7c330ef910_0 .net "out", 0 0, L_0x5c7c331614e0;  alias, 1 drivers
S_0x5c7c330effb0 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330ed4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330f0ff0_0 .net "in_a", 0 0, L_0x5c7c33161270;  alias, 1 drivers
v0x5c7c330f10c0_0 .net "in_b", 0 0, L_0x5c7c33161590;  alias, 1 drivers
v0x5c7c330f1190_0 .net "out", 0 0, L_0x5c7c33161800;  alias, 1 drivers
v0x5c7c330f12b0_0 .net "temp_out", 0 0, L_0x5c7c33161750;  1 drivers
S_0x5c7c330f0190 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330effb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161750 .functor NAND 1, L_0x5c7c33161270, L_0x5c7c33161590, C4<1>, C4<1>;
v0x5c7c330f03e0_0 .net "in_a", 0 0, L_0x5c7c33161270;  alias, 1 drivers
v0x5c7c330f04c0_0 .net "in_b", 0 0, L_0x5c7c33161590;  alias, 1 drivers
v0x5c7c330f0580_0 .net "out", 0 0, L_0x5c7c33161750;  alias, 1 drivers
S_0x5c7c330f06d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330effb0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f0e40_0 .net "in_a", 0 0, L_0x5c7c33161750;  alias, 1 drivers
v0x5c7c330f0ee0_0 .net "out", 0 0, L_0x5c7c33161800;  alias, 1 drivers
S_0x5c7c330f08f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f06d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161800 .functor NAND 1, L_0x5c7c33161750, L_0x5c7c33161750, C4<1>, C4<1>;
v0x5c7c330f0b60_0 .net "in_a", 0 0, L_0x5c7c33161750;  alias, 1 drivers
v0x5c7c330f0c50_0 .net "in_b", 0 0, L_0x5c7c33161750;  alias, 1 drivers
v0x5c7c330f0d40_0 .net "out", 0 0, L_0x5c7c33161800;  alias, 1 drivers
S_0x5c7c330f1400 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330ed4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f1b30_0 .net "in_a", 0 0, L_0x5c7c331611c0;  alias, 1 drivers
v0x5c7c330f1bd0_0 .net "out", 0 0, L_0x5c7c33161270;  alias, 1 drivers
S_0x5c7c330f15d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f1400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161270 .functor NAND 1, L_0x5c7c331611c0, L_0x5c7c331611c0, C4<1>, C4<1>;
v0x5c7c330f1840_0 .net "in_a", 0 0, L_0x5c7c331611c0;  alias, 1 drivers
v0x5c7c330f1900_0 .net "in_b", 0 0, L_0x5c7c331611c0;  alias, 1 drivers
v0x5c7c330f1a50_0 .net "out", 0 0, L_0x5c7c33161270;  alias, 1 drivers
S_0x5c7c330f1cd0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330ed4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f24a0_0 .net "in_a", 0 0, L_0x5c7c331614e0;  alias, 1 drivers
v0x5c7c330f2540_0 .net "out", 0 0, L_0x5c7c33161590;  alias, 1 drivers
S_0x5c7c330f1f40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f1cd0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161590 .functor NAND 1, L_0x5c7c331614e0, L_0x5c7c331614e0, C4<1>, C4<1>;
v0x5c7c330f21b0_0 .net "in_a", 0 0, L_0x5c7c331614e0;  alias, 1 drivers
v0x5c7c330f2270_0 .net "in_b", 0 0, L_0x5c7c331614e0;  alias, 1 drivers
v0x5c7c330f23c0_0 .net "out", 0 0, L_0x5c7c33161590;  alias, 1 drivers
S_0x5c7c330f2640 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330ed4b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f2de0_0 .net "in_a", 0 0, L_0x5c7c33161800;  alias, 1 drivers
v0x5c7c330f2e80_0 .net "out", 0 0, L_0x5c7c331618b0;  alias, 1 drivers
S_0x5c7c330f2860 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f2640;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331618b0 .functor NAND 1, L_0x5c7c33161800, L_0x5c7c33161800, C4<1>, C4<1>;
v0x5c7c330f2ad0_0 .net "in_a", 0 0, L_0x5c7c33161800;  alias, 1 drivers
v0x5c7c330f2b90_0 .net "in_b", 0 0, L_0x5c7c33161800;  alias, 1 drivers
v0x5c7c330f2ce0_0 .net "out", 0 0, L_0x5c7c331618b0;  alias, 1 drivers
S_0x5c7c330f3e20 .scope module, "mux_gate7" "Mux" 15 14, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c330fd180_0 .net "in_a", 0 0, L_0x5c7c33162890;  1 drivers
v0x5c7c330fd220_0 .net "in_b", 0 0, L_0x5c7c33162930;  1 drivers
v0x5c7c330fd330_0 .net "out", 0 0, L_0x5c7c331626d0;  1 drivers
v0x5c7c330fd3d0_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330fd470_0 .net "sel_out", 0 0, L_0x5c7c33160d30;  1 drivers
v0x5c7c330fd5f0_0 .net "temp_a_out", 0 0, L_0x5c7c33161d20;  1 drivers
v0x5c7c330fd7a0_0 .net "temp_b_out", 0 0, L_0x5c7c33161e80;  1 drivers
S_0x5c7c330f4020 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330f3e20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330f5080_0 .net "in_a", 0 0, L_0x5c7c33162890;  alias, 1 drivers
v0x5c7c330f5150_0 .net "in_b", 0 0, L_0x5c7c33160d30;  alias, 1 drivers
v0x5c7c330f5220_0 .net "out", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
v0x5c7c330f5340_0 .net "temp_out", 0 0, L_0x5c7c33161c70;  1 drivers
S_0x5c7c330f4290 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330f4020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161c70 .functor NAND 1, L_0x5c7c33162890, L_0x5c7c33160d30, C4<1>, C4<1>;
v0x5c7c330f4500_0 .net "in_a", 0 0, L_0x5c7c33162890;  alias, 1 drivers
v0x5c7c330f45e0_0 .net "in_b", 0 0, L_0x5c7c33160d30;  alias, 1 drivers
v0x5c7c330f46a0_0 .net "out", 0 0, L_0x5c7c33161c70;  alias, 1 drivers
S_0x5c7c330f47c0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330f4020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f4f00_0 .net "in_a", 0 0, L_0x5c7c33161c70;  alias, 1 drivers
v0x5c7c330f4fa0_0 .net "out", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
S_0x5c7c330f49e0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f47c0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161d20 .functor NAND 1, L_0x5c7c33161c70, L_0x5c7c33161c70, C4<1>, C4<1>;
v0x5c7c330f4c50_0 .net "in_a", 0 0, L_0x5c7c33161c70;  alias, 1 drivers
v0x5c7c330f4d10_0 .net "in_b", 0 0, L_0x5c7c33161c70;  alias, 1 drivers
v0x5c7c330f4e00_0 .net "out", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
S_0x5c7c330f5400 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330f3e20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330f6410_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330f64b0_0 .net "in_b", 0 0, L_0x5c7c33162930;  alias, 1 drivers
v0x5c7c330f65a0_0 .net "out", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
v0x5c7c330f66c0_0 .net "temp_out", 0 0, L_0x5c7c33161dd0;  1 drivers
S_0x5c7c330f55e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330f5400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161dd0 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33162930, C4<1>, C4<1>;
v0x5c7c330f5850_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330f5910_0 .net "in_b", 0 0, L_0x5c7c33162930;  alias, 1 drivers
v0x5c7c330f59d0_0 .net "out", 0 0, L_0x5c7c33161dd0;  alias, 1 drivers
S_0x5c7c330f5af0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330f5400;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f6260_0 .net "in_a", 0 0, L_0x5c7c33161dd0;  alias, 1 drivers
v0x5c7c330f6300_0 .net "out", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
S_0x5c7c330f5d10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f5af0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161e80 .functor NAND 1, L_0x5c7c33161dd0, L_0x5c7c33161dd0, C4<1>, C4<1>;
v0x5c7c330f5f80_0 .net "in_a", 0 0, L_0x5c7c33161dd0;  alias, 1 drivers
v0x5c7c330f6070_0 .net "in_b", 0 0, L_0x5c7c33161dd0;  alias, 1 drivers
v0x5c7c330f6160_0 .net "out", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
S_0x5c7c330f6780 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330f3e20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f6e80_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330f6f20_0 .net "out", 0 0, L_0x5c7c33160d30;  alias, 1 drivers
S_0x5c7c330f6950 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f6780;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33160d30 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c330f6ba0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330f6c60_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330f6d20_0 .net "out", 0 0, L_0x5c7c33160d30;  alias, 1 drivers
S_0x5c7c330f7020 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330f3e20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330fcad0_0 .net "branch1_out", 0 0, L_0x5c7c33162090;  1 drivers
v0x5c7c330fcc00_0 .net "branch2_out", 0 0, L_0x5c7c331623b0;  1 drivers
v0x5c7c330fcd50_0 .net "in_a", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
v0x5c7c330fce20_0 .net "in_b", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
v0x5c7c330fcec0_0 .net "out", 0 0, L_0x5c7c331626d0;  alias, 1 drivers
v0x5c7c330fcf60_0 .net "temp1_out", 0 0, L_0x5c7c33161fe0;  1 drivers
v0x5c7c330fd000_0 .net "temp2_out", 0 0, L_0x5c7c33162300;  1 drivers
v0x5c7c330fd0a0_0 .net "temp3_out", 0 0, L_0x5c7c33162620;  1 drivers
S_0x5c7c330f7250 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c330f7020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330f8310_0 .net "in_a", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
v0x5c7c330f83b0_0 .net "in_b", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
v0x5c7c330f8470_0 .net "out", 0 0, L_0x5c7c33161fe0;  alias, 1 drivers
v0x5c7c330f8590_0 .net "temp_out", 0 0, L_0x5c7c33161f30;  1 drivers
S_0x5c7c330f74c0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330f7250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161f30 .functor NAND 1, L_0x5c7c33161d20, L_0x5c7c33161d20, C4<1>, C4<1>;
v0x5c7c330f7730_0 .net "in_a", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
v0x5c7c330f77f0_0 .net "in_b", 0 0, L_0x5c7c33161d20;  alias, 1 drivers
v0x5c7c330f7940_0 .net "out", 0 0, L_0x5c7c33161f30;  alias, 1 drivers
S_0x5c7c330f7a40 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330f7250;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f8160_0 .net "in_a", 0 0, L_0x5c7c33161f30;  alias, 1 drivers
v0x5c7c330f8200_0 .net "out", 0 0, L_0x5c7c33161fe0;  alias, 1 drivers
S_0x5c7c330f7c10 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f7a40;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33161fe0 .functor NAND 1, L_0x5c7c33161f30, L_0x5c7c33161f30, C4<1>, C4<1>;
v0x5c7c330f7e80_0 .net "in_a", 0 0, L_0x5c7c33161f30;  alias, 1 drivers
v0x5c7c330f7f70_0 .net "in_b", 0 0, L_0x5c7c33161f30;  alias, 1 drivers
v0x5c7c330f8060_0 .net "out", 0 0, L_0x5c7c33161fe0;  alias, 1 drivers
S_0x5c7c330f8700 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c330f7020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330f9730_0 .net "in_a", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
v0x5c7c330f97d0_0 .net "in_b", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
v0x5c7c330f9890_0 .net "out", 0 0, L_0x5c7c33162300;  alias, 1 drivers
v0x5c7c330f99b0_0 .net "temp_out", 0 0, L_0x5c7c33162250;  1 drivers
S_0x5c7c330f88e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330f8700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162250 .functor NAND 1, L_0x5c7c33161e80, L_0x5c7c33161e80, C4<1>, C4<1>;
v0x5c7c330f8b50_0 .net "in_a", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
v0x5c7c330f8c10_0 .net "in_b", 0 0, L_0x5c7c33161e80;  alias, 1 drivers
v0x5c7c330f8d60_0 .net "out", 0 0, L_0x5c7c33162250;  alias, 1 drivers
S_0x5c7c330f8e60 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330f8700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330f9580_0 .net "in_a", 0 0, L_0x5c7c33162250;  alias, 1 drivers
v0x5c7c330f9620_0 .net "out", 0 0, L_0x5c7c33162300;  alias, 1 drivers
S_0x5c7c330f9030 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330f8e60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162300 .functor NAND 1, L_0x5c7c33162250, L_0x5c7c33162250, C4<1>, C4<1>;
v0x5c7c330f92a0_0 .net "in_a", 0 0, L_0x5c7c33162250;  alias, 1 drivers
v0x5c7c330f9390_0 .net "in_b", 0 0, L_0x5c7c33162250;  alias, 1 drivers
v0x5c7c330f9480_0 .net "out", 0 0, L_0x5c7c33162300;  alias, 1 drivers
S_0x5c7c330f9b20 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c330f7020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330fab60_0 .net "in_a", 0 0, L_0x5c7c33162090;  alias, 1 drivers
v0x5c7c330fac30_0 .net "in_b", 0 0, L_0x5c7c331623b0;  alias, 1 drivers
v0x5c7c330fad00_0 .net "out", 0 0, L_0x5c7c33162620;  alias, 1 drivers
v0x5c7c330fae20_0 .net "temp_out", 0 0, L_0x5c7c33162570;  1 drivers
S_0x5c7c330f9d00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330f9b20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162570 .functor NAND 1, L_0x5c7c33162090, L_0x5c7c331623b0, C4<1>, C4<1>;
v0x5c7c330f9f50_0 .net "in_a", 0 0, L_0x5c7c33162090;  alias, 1 drivers
v0x5c7c330fa030_0 .net "in_b", 0 0, L_0x5c7c331623b0;  alias, 1 drivers
v0x5c7c330fa0f0_0 .net "out", 0 0, L_0x5c7c33162570;  alias, 1 drivers
S_0x5c7c330fa240 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330f9b20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330fa9b0_0 .net "in_a", 0 0, L_0x5c7c33162570;  alias, 1 drivers
v0x5c7c330faa50_0 .net "out", 0 0, L_0x5c7c33162620;  alias, 1 drivers
S_0x5c7c330fa460 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330fa240;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162620 .functor NAND 1, L_0x5c7c33162570, L_0x5c7c33162570, C4<1>, C4<1>;
v0x5c7c330fa6d0_0 .net "in_a", 0 0, L_0x5c7c33162570;  alias, 1 drivers
v0x5c7c330fa7c0_0 .net "in_b", 0 0, L_0x5c7c33162570;  alias, 1 drivers
v0x5c7c330fa8b0_0 .net "out", 0 0, L_0x5c7c33162620;  alias, 1 drivers
S_0x5c7c330faf70 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c330f7020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330fb6a0_0 .net "in_a", 0 0, L_0x5c7c33161fe0;  alias, 1 drivers
v0x5c7c330fb740_0 .net "out", 0 0, L_0x5c7c33162090;  alias, 1 drivers
S_0x5c7c330fb140 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330faf70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162090 .functor NAND 1, L_0x5c7c33161fe0, L_0x5c7c33161fe0, C4<1>, C4<1>;
v0x5c7c330fb3b0_0 .net "in_a", 0 0, L_0x5c7c33161fe0;  alias, 1 drivers
v0x5c7c330fb470_0 .net "in_b", 0 0, L_0x5c7c33161fe0;  alias, 1 drivers
v0x5c7c330fb5c0_0 .net "out", 0 0, L_0x5c7c33162090;  alias, 1 drivers
S_0x5c7c330fb840 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c330f7020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330fc010_0 .net "in_a", 0 0, L_0x5c7c33162300;  alias, 1 drivers
v0x5c7c330fc0b0_0 .net "out", 0 0, L_0x5c7c331623b0;  alias, 1 drivers
S_0x5c7c330fbab0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330fb840;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331623b0 .functor NAND 1, L_0x5c7c33162300, L_0x5c7c33162300, C4<1>, C4<1>;
v0x5c7c330fbd20_0 .net "in_a", 0 0, L_0x5c7c33162300;  alias, 1 drivers
v0x5c7c330fbde0_0 .net "in_b", 0 0, L_0x5c7c33162300;  alias, 1 drivers
v0x5c7c330fbf30_0 .net "out", 0 0, L_0x5c7c331623b0;  alias, 1 drivers
S_0x5c7c330fc1b0 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c330f7020;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330fc950_0 .net "in_a", 0 0, L_0x5c7c33162620;  alias, 1 drivers
v0x5c7c330fc9f0_0 .net "out", 0 0, L_0x5c7c331626d0;  alias, 1 drivers
S_0x5c7c330fc3d0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330fc1b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331626d0 .functor NAND 1, L_0x5c7c33162620, L_0x5c7c33162620, C4<1>, C4<1>;
v0x5c7c330fc640_0 .net "in_a", 0 0, L_0x5c7c33162620;  alias, 1 drivers
v0x5c7c330fc700_0 .net "in_b", 0 0, L_0x5c7c33162620;  alias, 1 drivers
v0x5c7c330fc850_0 .net "out", 0 0, L_0x5c7c331626d0;  alias, 1 drivers
S_0x5c7c330fd990 .scope module, "mux_gate8" "Mux" 15 15, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33106cf0_0 .net "in_a", 0 0, L_0x5c7c33163730;  1 drivers
v0x5c7c33106d90_0 .net "in_b", 0 0, L_0x5c7c331637d0;  1 drivers
v0x5c7c33106ea0_0 .net "out", 0 0, L_0x5c7c33163570;  1 drivers
v0x5c7c33106f40_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33106fe0_0 .net "sel_out", 0 0, L_0x5c7c33162a60;  1 drivers
v0x5c7c33107160_0 .net "temp_a_out", 0 0, L_0x5c7c33162bc0;  1 drivers
v0x5c7c33107310_0 .net "temp_b_out", 0 0, L_0x5c7c33162d20;  1 drivers
S_0x5c7c330fdb90 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c330fd990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330febf0_0 .net "in_a", 0 0, L_0x5c7c33163730;  alias, 1 drivers
v0x5c7c330fecc0_0 .net "in_b", 0 0, L_0x5c7c33162a60;  alias, 1 drivers
v0x5c7c330fed90_0 .net "out", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
v0x5c7c330feeb0_0 .net "temp_out", 0 0, L_0x5c7c33162b10;  1 drivers
S_0x5c7c330fde00 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330fdb90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162b10 .functor NAND 1, L_0x5c7c33163730, L_0x5c7c33162a60, C4<1>, C4<1>;
v0x5c7c330fe070_0 .net "in_a", 0 0, L_0x5c7c33163730;  alias, 1 drivers
v0x5c7c330fe150_0 .net "in_b", 0 0, L_0x5c7c33162a60;  alias, 1 drivers
v0x5c7c330fe210_0 .net "out", 0 0, L_0x5c7c33162b10;  alias, 1 drivers
S_0x5c7c330fe330 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330fdb90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330fea70_0 .net "in_a", 0 0, L_0x5c7c33162b10;  alias, 1 drivers
v0x5c7c330feb10_0 .net "out", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
S_0x5c7c330fe550 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330fe330;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162bc0 .functor NAND 1, L_0x5c7c33162b10, L_0x5c7c33162b10, C4<1>, C4<1>;
v0x5c7c330fe7c0_0 .net "in_a", 0 0, L_0x5c7c33162b10;  alias, 1 drivers
v0x5c7c330fe880_0 .net "in_b", 0 0, L_0x5c7c33162b10;  alias, 1 drivers
v0x5c7c330fe970_0 .net "out", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
S_0x5c7c330fef70 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c330fd990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c330fff80_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33100020_0 .net "in_b", 0 0, L_0x5c7c331637d0;  alias, 1 drivers
v0x5c7c33100110_0 .net "out", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
v0x5c7c33100230_0 .net "temp_out", 0 0, L_0x5c7c33162c70;  1 drivers
S_0x5c7c330ff150 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c330fef70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162c70 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c331637d0, C4<1>, C4<1>;
v0x5c7c330ff3c0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c330ff480_0 .net "in_b", 0 0, L_0x5c7c331637d0;  alias, 1 drivers
v0x5c7c330ff540_0 .net "out", 0 0, L_0x5c7c33162c70;  alias, 1 drivers
S_0x5c7c330ff660 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c330fef70;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c330ffdd0_0 .net "in_a", 0 0, L_0x5c7c33162c70;  alias, 1 drivers
v0x5c7c330ffe70_0 .net "out", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
S_0x5c7c330ff880 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c330ff660;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162d20 .functor NAND 1, L_0x5c7c33162c70, L_0x5c7c33162c70, C4<1>, C4<1>;
v0x5c7c330ffaf0_0 .net "in_a", 0 0, L_0x5c7c33162c70;  alias, 1 drivers
v0x5c7c330ffbe0_0 .net "in_b", 0 0, L_0x5c7c33162c70;  alias, 1 drivers
v0x5c7c330ffcd0_0 .net "out", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
S_0x5c7c331002f0 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c330fd990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c331009f0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33100a90_0 .net "out", 0 0, L_0x5c7c33162a60;  alias, 1 drivers
S_0x5c7c331004c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c331002f0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162a60 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c33100710_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c331007d0_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33100890_0 .net "out", 0 0, L_0x5c7c33162a60;  alias, 1 drivers
S_0x5c7c33100b90 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c330fd990;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33106640_0 .net "branch1_out", 0 0, L_0x5c7c33162f30;  1 drivers
v0x5c7c33106770_0 .net "branch2_out", 0 0, L_0x5c7c33163250;  1 drivers
v0x5c7c331068c0_0 .net "in_a", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
v0x5c7c33106990_0 .net "in_b", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
v0x5c7c33106a30_0 .net "out", 0 0, L_0x5c7c33163570;  alias, 1 drivers
v0x5c7c33106ad0_0 .net "temp1_out", 0 0, L_0x5c7c33162e80;  1 drivers
v0x5c7c33106b70_0 .net "temp2_out", 0 0, L_0x5c7c331631a0;  1 drivers
v0x5c7c33106c10_0 .net "temp3_out", 0 0, L_0x5c7c331634c0;  1 drivers
S_0x5c7c33100dc0 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c33100b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33101e80_0 .net "in_a", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
v0x5c7c33101f20_0 .net "in_b", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
v0x5c7c33101fe0_0 .net "out", 0 0, L_0x5c7c33162e80;  alias, 1 drivers
v0x5c7c33102100_0 .net "temp_out", 0 0, L_0x5c7c33162dd0;  1 drivers
S_0x5c7c33101030 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33100dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162dd0 .functor NAND 1, L_0x5c7c33162bc0, L_0x5c7c33162bc0, C4<1>, C4<1>;
v0x5c7c331012a0_0 .net "in_a", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
v0x5c7c33101360_0 .net "in_b", 0 0, L_0x5c7c33162bc0;  alias, 1 drivers
v0x5c7c331014b0_0 .net "out", 0 0, L_0x5c7c33162dd0;  alias, 1 drivers
S_0x5c7c331015b0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33100dc0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33101cd0_0 .net "in_a", 0 0, L_0x5c7c33162dd0;  alias, 1 drivers
v0x5c7c33101d70_0 .net "out", 0 0, L_0x5c7c33162e80;  alias, 1 drivers
S_0x5c7c33101780 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c331015b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162e80 .functor NAND 1, L_0x5c7c33162dd0, L_0x5c7c33162dd0, C4<1>, C4<1>;
v0x5c7c331019f0_0 .net "in_a", 0 0, L_0x5c7c33162dd0;  alias, 1 drivers
v0x5c7c33101ae0_0 .net "in_b", 0 0, L_0x5c7c33162dd0;  alias, 1 drivers
v0x5c7c33101bd0_0 .net "out", 0 0, L_0x5c7c33162e80;  alias, 1 drivers
S_0x5c7c33102270 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c33100b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c331032a0_0 .net "in_a", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
v0x5c7c33103340_0 .net "in_b", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
v0x5c7c33103400_0 .net "out", 0 0, L_0x5c7c331631a0;  alias, 1 drivers
v0x5c7c33103520_0 .net "temp_out", 0 0, L_0x5c7c331630f0;  1 drivers
S_0x5c7c33102450 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33102270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331630f0 .functor NAND 1, L_0x5c7c33162d20, L_0x5c7c33162d20, C4<1>, C4<1>;
v0x5c7c331026c0_0 .net "in_a", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
v0x5c7c33102780_0 .net "in_b", 0 0, L_0x5c7c33162d20;  alias, 1 drivers
v0x5c7c331028d0_0 .net "out", 0 0, L_0x5c7c331630f0;  alias, 1 drivers
S_0x5c7c331029d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33102270;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c331030f0_0 .net "in_a", 0 0, L_0x5c7c331630f0;  alias, 1 drivers
v0x5c7c33103190_0 .net "out", 0 0, L_0x5c7c331631a0;  alias, 1 drivers
S_0x5c7c33102ba0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c331029d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331631a0 .functor NAND 1, L_0x5c7c331630f0, L_0x5c7c331630f0, C4<1>, C4<1>;
v0x5c7c33102e10_0 .net "in_a", 0 0, L_0x5c7c331630f0;  alias, 1 drivers
v0x5c7c33102f00_0 .net "in_b", 0 0, L_0x5c7c331630f0;  alias, 1 drivers
v0x5c7c33102ff0_0 .net "out", 0 0, L_0x5c7c331631a0;  alias, 1 drivers
S_0x5c7c33103690 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c33100b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c331046d0_0 .net "in_a", 0 0, L_0x5c7c33162f30;  alias, 1 drivers
v0x5c7c331047a0_0 .net "in_b", 0 0, L_0x5c7c33163250;  alias, 1 drivers
v0x5c7c33104870_0 .net "out", 0 0, L_0x5c7c331634c0;  alias, 1 drivers
v0x5c7c33104990_0 .net "temp_out", 0 0, L_0x5c7c33163410;  1 drivers
S_0x5c7c33103870 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33103690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163410 .functor NAND 1, L_0x5c7c33162f30, L_0x5c7c33163250, C4<1>, C4<1>;
v0x5c7c33103ac0_0 .net "in_a", 0 0, L_0x5c7c33162f30;  alias, 1 drivers
v0x5c7c33103ba0_0 .net "in_b", 0 0, L_0x5c7c33163250;  alias, 1 drivers
v0x5c7c33103c60_0 .net "out", 0 0, L_0x5c7c33163410;  alias, 1 drivers
S_0x5c7c33103db0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33103690;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33104520_0 .net "in_a", 0 0, L_0x5c7c33163410;  alias, 1 drivers
v0x5c7c331045c0_0 .net "out", 0 0, L_0x5c7c331634c0;  alias, 1 drivers
S_0x5c7c33103fd0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33103db0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331634c0 .functor NAND 1, L_0x5c7c33163410, L_0x5c7c33163410, C4<1>, C4<1>;
v0x5c7c33104240_0 .net "in_a", 0 0, L_0x5c7c33163410;  alias, 1 drivers
v0x5c7c33104330_0 .net "in_b", 0 0, L_0x5c7c33163410;  alias, 1 drivers
v0x5c7c33104420_0 .net "out", 0 0, L_0x5c7c331634c0;  alias, 1 drivers
S_0x5c7c33104ae0 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c33100b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33105210_0 .net "in_a", 0 0, L_0x5c7c33162e80;  alias, 1 drivers
v0x5c7c331052b0_0 .net "out", 0 0, L_0x5c7c33162f30;  alias, 1 drivers
S_0x5c7c33104cb0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33104ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33162f30 .functor NAND 1, L_0x5c7c33162e80, L_0x5c7c33162e80, C4<1>, C4<1>;
v0x5c7c33104f20_0 .net "in_a", 0 0, L_0x5c7c33162e80;  alias, 1 drivers
v0x5c7c33104fe0_0 .net "in_b", 0 0, L_0x5c7c33162e80;  alias, 1 drivers
v0x5c7c33105130_0 .net "out", 0 0, L_0x5c7c33162f30;  alias, 1 drivers
S_0x5c7c331053b0 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c33100b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33105b80_0 .net "in_a", 0 0, L_0x5c7c331631a0;  alias, 1 drivers
v0x5c7c33105c20_0 .net "out", 0 0, L_0x5c7c33163250;  alias, 1 drivers
S_0x5c7c33105620 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c331053b0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163250 .functor NAND 1, L_0x5c7c331631a0, L_0x5c7c331631a0, C4<1>, C4<1>;
v0x5c7c33105890_0 .net "in_a", 0 0, L_0x5c7c331631a0;  alias, 1 drivers
v0x5c7c33105950_0 .net "in_b", 0 0, L_0x5c7c331631a0;  alias, 1 drivers
v0x5c7c33105aa0_0 .net "out", 0 0, L_0x5c7c33163250;  alias, 1 drivers
S_0x5c7c33105d20 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c33100b90;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c331064c0_0 .net "in_a", 0 0, L_0x5c7c331634c0;  alias, 1 drivers
v0x5c7c33106560_0 .net "out", 0 0, L_0x5c7c33163570;  alias, 1 drivers
S_0x5c7c33105f40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33105d20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163570 .functor NAND 1, L_0x5c7c331634c0, L_0x5c7c331634c0, C4<1>, C4<1>;
v0x5c7c331061b0_0 .net "in_a", 0 0, L_0x5c7c331634c0;  alias, 1 drivers
v0x5c7c33106270_0 .net "in_b", 0 0, L_0x5c7c331634c0;  alias, 1 drivers
v0x5c7c331063c0_0 .net "out", 0 0, L_0x5c7c33163570;  alias, 1 drivers
S_0x5c7c33107500 .scope module, "mux_gate9" "Mux" 15 16, 16 3 0, S_0x5c7c33054df0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
    .port_info 3 /INPUT 1 "sel";
v0x5c7c33110860_0 .net "in_a", 0 0, L_0x5c7c331645e0;  1 drivers
v0x5c7c33110900_0 .net "in_b", 0 0, L_0x5c7c33164680;  1 drivers
v0x5c7c33110a10_0 .net "out", 0 0, L_0x5c7c33164420;  1 drivers
v0x5c7c33110ab0_0 .net "sel", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33110b50_0 .net "sel_out", 0 0, L_0x5c7c33163910;  1 drivers
v0x5c7c33110cd0_0 .net "temp_a_out", 0 0, L_0x5c7c33163a70;  1 drivers
v0x5c7c33110e80_0 .net "temp_b_out", 0 0, L_0x5c7c33163bd0;  1 drivers
S_0x5c7c33107700 .scope module, "and_gate" "And" 16 9, 5 2 0, S_0x5c7c33107500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33108760_0 .net "in_a", 0 0, L_0x5c7c331645e0;  alias, 1 drivers
v0x5c7c33108830_0 .net "in_b", 0 0, L_0x5c7c33163910;  alias, 1 drivers
v0x5c7c33108900_0 .net "out", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
v0x5c7c33108a20_0 .net "temp_out", 0 0, L_0x5c7c331639c0;  1 drivers
S_0x5c7c33107970 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33107700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331639c0 .functor NAND 1, L_0x5c7c331645e0, L_0x5c7c33163910, C4<1>, C4<1>;
v0x5c7c33107be0_0 .net "in_a", 0 0, L_0x5c7c331645e0;  alias, 1 drivers
v0x5c7c33107cc0_0 .net "in_b", 0 0, L_0x5c7c33163910;  alias, 1 drivers
v0x5c7c33107d80_0 .net "out", 0 0, L_0x5c7c331639c0;  alias, 1 drivers
S_0x5c7c33107ea0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33107700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c331085e0_0 .net "in_a", 0 0, L_0x5c7c331639c0;  alias, 1 drivers
v0x5c7c33108680_0 .net "out", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
S_0x5c7c331080c0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33107ea0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163a70 .functor NAND 1, L_0x5c7c331639c0, L_0x5c7c331639c0, C4<1>, C4<1>;
v0x5c7c33108330_0 .net "in_a", 0 0, L_0x5c7c331639c0;  alias, 1 drivers
v0x5c7c331083f0_0 .net "in_b", 0 0, L_0x5c7c331639c0;  alias, 1 drivers
v0x5c7c331084e0_0 .net "out", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
S_0x5c7c33108ae0 .scope module, "and_gate3" "And" 16 10, 5 2 0, S_0x5c7c33107500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c33109af0_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33109b90_0 .net "in_b", 0 0, L_0x5c7c33164680;  alias, 1 drivers
v0x5c7c33109c80_0 .net "out", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
v0x5c7c33109da0_0 .net "temp_out", 0 0, L_0x5c7c33163b20;  1 drivers
S_0x5c7c33108cc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c33108ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163b20 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33164680, C4<1>, C4<1>;
v0x5c7c33108f30_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c33108ff0_0 .net "in_b", 0 0, L_0x5c7c33164680;  alias, 1 drivers
v0x5c7c331090b0_0 .net "out", 0 0, L_0x5c7c33163b20;  alias, 1 drivers
S_0x5c7c331091d0 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c33108ae0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33109940_0 .net "in_a", 0 0, L_0x5c7c33163b20;  alias, 1 drivers
v0x5c7c331099e0_0 .net "out", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
S_0x5c7c331093f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c331091d0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163bd0 .functor NAND 1, L_0x5c7c33163b20, L_0x5c7c33163b20, C4<1>, C4<1>;
v0x5c7c33109660_0 .net "in_a", 0 0, L_0x5c7c33163b20;  alias, 1 drivers
v0x5c7c33109750_0 .net "in_b", 0 0, L_0x5c7c33163b20;  alias, 1 drivers
v0x5c7c33109840_0 .net "out", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
S_0x5c7c33109e60 .scope module, "not_gate2" "Not" 16 8, 7 3 0, S_0x5c7c33107500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3310a560_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3310a600_0 .net "out", 0 0, L_0x5c7c33163910;  alias, 1 drivers
S_0x5c7c3310a030 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c33109e60;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163910 .functor NAND 1, L_0x5c7c33169ff0, L_0x5c7c33169ff0, C4<1>, C4<1>;
v0x5c7c3310a280_0 .net "in_a", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3310a340_0 .net "in_b", 0 0, L_0x5c7c33169ff0;  alias, 1 drivers
v0x5c7c3310a400_0 .net "out", 0 0, L_0x5c7c33163910;  alias, 1 drivers
S_0x5c7c3310a700 .scope module, "or_gate" "Or" 16 11, 9 3 0, S_0x5c7c33107500;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c331101b0_0 .net "branch1_out", 0 0, L_0x5c7c33163de0;  1 drivers
v0x5c7c331102e0_0 .net "branch2_out", 0 0, L_0x5c7c33164100;  1 drivers
v0x5c7c33110430_0 .net "in_a", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
v0x5c7c33110500_0 .net "in_b", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
v0x5c7c331105a0_0 .net "out", 0 0, L_0x5c7c33164420;  alias, 1 drivers
v0x5c7c33110640_0 .net "temp1_out", 0 0, L_0x5c7c33163d30;  1 drivers
v0x5c7c331106e0_0 .net "temp2_out", 0 0, L_0x5c7c33164050;  1 drivers
v0x5c7c33110780_0 .net "temp3_out", 0 0, L_0x5c7c33164370;  1 drivers
S_0x5c7c3310a930 .scope module, "and_gate" "And" 9 9, 5 2 0, S_0x5c7c3310a700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3310b9f0_0 .net "in_a", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
v0x5c7c3310ba90_0 .net "in_b", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
v0x5c7c3310bb50_0 .net "out", 0 0, L_0x5c7c33163d30;  alias, 1 drivers
v0x5c7c3310bc70_0 .net "temp_out", 0 0, L_0x5c7c33163c80;  1 drivers
S_0x5c7c3310aba0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3310a930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163c80 .functor NAND 1, L_0x5c7c33163a70, L_0x5c7c33163a70, C4<1>, C4<1>;
v0x5c7c3310ae10_0 .net "in_a", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
v0x5c7c3310aed0_0 .net "in_b", 0 0, L_0x5c7c33163a70;  alias, 1 drivers
v0x5c7c3310b020_0 .net "out", 0 0, L_0x5c7c33163c80;  alias, 1 drivers
S_0x5c7c3310b120 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3310a930;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3310b840_0 .net "in_a", 0 0, L_0x5c7c33163c80;  alias, 1 drivers
v0x5c7c3310b8e0_0 .net "out", 0 0, L_0x5c7c33163d30;  alias, 1 drivers
S_0x5c7c3310b2f0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3310b120;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163d30 .functor NAND 1, L_0x5c7c33163c80, L_0x5c7c33163c80, C4<1>, C4<1>;
v0x5c7c3310b560_0 .net "in_a", 0 0, L_0x5c7c33163c80;  alias, 1 drivers
v0x5c7c3310b650_0 .net "in_b", 0 0, L_0x5c7c33163c80;  alias, 1 drivers
v0x5c7c3310b740_0 .net "out", 0 0, L_0x5c7c33163d30;  alias, 1 drivers
S_0x5c7c3310bde0 .scope module, "and_gate2" "And" 9 13, 5 2 0, S_0x5c7c3310a700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3310ce10_0 .net "in_a", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
v0x5c7c3310ceb0_0 .net "in_b", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
v0x5c7c3310cf70_0 .net "out", 0 0, L_0x5c7c33164050;  alias, 1 drivers
v0x5c7c3310d090_0 .net "temp_out", 0 0, L_0x5c7c33163fa0;  1 drivers
S_0x5c7c3310bfc0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3310bde0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163fa0 .functor NAND 1, L_0x5c7c33163bd0, L_0x5c7c33163bd0, C4<1>, C4<1>;
v0x5c7c3310c230_0 .net "in_a", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
v0x5c7c3310c2f0_0 .net "in_b", 0 0, L_0x5c7c33163bd0;  alias, 1 drivers
v0x5c7c3310c440_0 .net "out", 0 0, L_0x5c7c33163fa0;  alias, 1 drivers
S_0x5c7c3310c540 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3310bde0;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3310cc60_0 .net "in_a", 0 0, L_0x5c7c33163fa0;  alias, 1 drivers
v0x5c7c3310cd00_0 .net "out", 0 0, L_0x5c7c33164050;  alias, 1 drivers
S_0x5c7c3310c710 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3310c540;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33164050 .functor NAND 1, L_0x5c7c33163fa0, L_0x5c7c33163fa0, C4<1>, C4<1>;
v0x5c7c3310c980_0 .net "in_a", 0 0, L_0x5c7c33163fa0;  alias, 1 drivers
v0x5c7c3310ca70_0 .net "in_b", 0 0, L_0x5c7c33163fa0;  alias, 1 drivers
v0x5c7c3310cb60_0 .net "out", 0 0, L_0x5c7c33164050;  alias, 1 drivers
S_0x5c7c3310d200 .scope module, "and_gate3" "And" 9 17, 5 2 0, S_0x5c7c3310a700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
v0x5c7c3310e240_0 .net "in_a", 0 0, L_0x5c7c33163de0;  alias, 1 drivers
v0x5c7c3310e310_0 .net "in_b", 0 0, L_0x5c7c33164100;  alias, 1 drivers
v0x5c7c3310e3e0_0 .net "out", 0 0, L_0x5c7c33164370;  alias, 1 drivers
v0x5c7c3310e500_0 .net "temp_out", 0 0, L_0x5c7c331642c0;  1 drivers
S_0x5c7c3310d3e0 .scope module, "nand_gate" "Nand" 5 7, 6 1 0, S_0x5c7c3310d200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c331642c0 .functor NAND 1, L_0x5c7c33163de0, L_0x5c7c33164100, C4<1>, C4<1>;
v0x5c7c3310d630_0 .net "in_a", 0 0, L_0x5c7c33163de0;  alias, 1 drivers
v0x5c7c3310d710_0 .net "in_b", 0 0, L_0x5c7c33164100;  alias, 1 drivers
v0x5c7c3310d7d0_0 .net "out", 0 0, L_0x5c7c331642c0;  alias, 1 drivers
S_0x5c7c3310d920 .scope module, "not_gate" "Not" 5 8, 7 3 0, S_0x5c7c3310d200;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3310e090_0 .net "in_a", 0 0, L_0x5c7c331642c0;  alias, 1 drivers
v0x5c7c3310e130_0 .net "out", 0 0, L_0x5c7c33164370;  alias, 1 drivers
S_0x5c7c3310db40 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3310d920;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33164370 .functor NAND 1, L_0x5c7c331642c0, L_0x5c7c331642c0, C4<1>, C4<1>;
v0x5c7c3310ddb0_0 .net "in_a", 0 0, L_0x5c7c331642c0;  alias, 1 drivers
v0x5c7c3310dea0_0 .net "in_b", 0 0, L_0x5c7c331642c0;  alias, 1 drivers
v0x5c7c3310df90_0 .net "out", 0 0, L_0x5c7c33164370;  alias, 1 drivers
S_0x5c7c3310e650 .scope module, "not_gate" "Not" 9 10, 7 3 0, S_0x5c7c3310a700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3310ed80_0 .net "in_a", 0 0, L_0x5c7c33163d30;  alias, 1 drivers
v0x5c7c3310ee20_0 .net "out", 0 0, L_0x5c7c33163de0;  alias, 1 drivers
S_0x5c7c3310e820 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3310e650;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33163de0 .functor NAND 1, L_0x5c7c33163d30, L_0x5c7c33163d30, C4<1>, C4<1>;
v0x5c7c3310ea90_0 .net "in_a", 0 0, L_0x5c7c33163d30;  alias, 1 drivers
v0x5c7c3310eb50_0 .net "in_b", 0 0, L_0x5c7c33163d30;  alias, 1 drivers
v0x5c7c3310eca0_0 .net "out", 0 0, L_0x5c7c33163de0;  alias, 1 drivers
S_0x5c7c3310ef20 .scope module, "not_gate2" "Not" 9 14, 7 3 0, S_0x5c7c3310a700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c3310f6f0_0 .net "in_a", 0 0, L_0x5c7c33164050;  alias, 1 drivers
v0x5c7c3310f790_0 .net "out", 0 0, L_0x5c7c33164100;  alias, 1 drivers
S_0x5c7c3310f190 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3310ef20;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33164100 .functor NAND 1, L_0x5c7c33164050, L_0x5c7c33164050, C4<1>, C4<1>;
v0x5c7c3310f400_0 .net "in_a", 0 0, L_0x5c7c33164050;  alias, 1 drivers
v0x5c7c3310f4c0_0 .net "in_b", 0 0, L_0x5c7c33164050;  alias, 1 drivers
v0x5c7c3310f610_0 .net "out", 0 0, L_0x5c7c33164100;  alias, 1 drivers
S_0x5c7c3310f890 .scope module, "not_gate3" "Not" 9 18, 7 3 0, S_0x5c7c3310a700;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /OUTPUT 1 "out";
v0x5c7c33110030_0 .net "in_a", 0 0, L_0x5c7c33164370;  alias, 1 drivers
v0x5c7c331100d0_0 .net "out", 0 0, L_0x5c7c33164420;  alias, 1 drivers
S_0x5c7c3310fab0 .scope module, "nand_gate" "Nand" 7 7, 6 1 0, S_0x5c7c3310f890;
 .timescale 0 0;
    .port_info 0 /INPUT 1 "in_a";
    .port_info 1 /INPUT 1 "in_b";
    .port_info 2 /OUTPUT 1 "out";
L_0x5c7c33164420 .functor NAND 1, L_0x5c7c33164370, L_0x5c7c33164370, C4<1>, C4<1>;
v0x5c7c3310fd20_0 .net "in_a", 0 0, L_0x5c7c33164370;  alias, 1 drivers
v0x5c7c3310fde0_0 .net "in_b", 0 0, L_0x5c7c33164370;  alias, 1 drivers
v0x5c7c3310ff30_0 .net "out", 0 0, L_0x5c7c33164420;  alias, 1 drivers
# The file index is used to find the file name in the following table.
:file_names 17;
    "N/A";
    "<interactive>";
    "./Add16/src/Add16.vh";
    "./FullAdder/src/FullAdder.vh";
    "./HalfAdder/src/HalfAdder.vh";
    "./And/src/And.vh";
    "./Nand/src/Nand.vh";
    "./Not/src/Not.vh";
    "./Xor/src/Xor.vh";
    "./Or/src/Or.vh";
    "./And16/src/And16.vh";
    "./Not16/src/Not16.vh";
    "./DMux4Way/src/DMux4Way.vh";
    "./DMux/src/DMux.vh";
    "./Mux4Way16/src/Mux4Way16.vh";
    "Mux16/src/Mux16.vh";
    "./Mux/src/Mux.vh";
