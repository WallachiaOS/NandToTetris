module Nand(in_a,in_b,out);
    input in_a,in_b;
    output out;
    
    nand(out,in_a,in_b);
endmodule